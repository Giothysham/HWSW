--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"004124230031222300112023340111730000001300000013000000131140006f",
        INIT_01 => X"02c1242302b1222302a1202300912e2300812c2300712a230061282300512623",
        INIT_02 => X"05412423053122230521202303112e2303012c2302f12a2302e1282302d12623",
        INIT_03 => X"07c1242307b1222307a1202305912e2305812c2305712a230561282305512623",
        INIT_04 => X"008122030041218300012083278000ef3420357307f12a2307e1282307d12623",
        INIT_05 => X"02812603024125830201250301c1248301812403014123830101230300c12283",
        INIT_06 => X"04812a03044129830401290303c1288303812803034127830301270302c12683",
        INIT_07 => X"06812e0306412d8306012d0305c12c8305812c0305412b8305012b0304c12a83",
        INIT_08 => X"000001930000011300000093302000733401117307412f8307012f0306c12e83",
        INIT_09 => X"0000059300000513000004930000041300000393000003130000029300000213",
        INIT_0A => X"0000099300000913000008930000081300000793000007130000069300000613",
        INIT_0B => X"00000d9300000d1300000c9300000c1300000b9300000b1300000a9300000a13",
        INIT_0C => X"0000113700018213eef18193deadc1b700000f9300000f1300000e9300000e13",
        INIT_0D => X"30411073fff001133004507330511073e6810113000001173401107300010113",
        INIT_0E => X"00112023ff4101130540006f7ac000ef001000737b4000effe01011300001137",
        INIT_0F => X"0005853300029663fff50293000583330280006f000514630061242300512223",
        INIT_10 => X"00812303004122830001208300030533fe029ce3fff2829300b303330140006f",
        INIT_11 => X"810007b70101041300812623ff0101130000006f0000006f0000806700c10113",
        INIT_12 => X"000080670101011300c124030000001300e7a02300776713810007b70007a703",
        INIT_13 => X"810007b70007a703810007b7068000ef010104130081242300112623ff010113",
        INIT_14 => X"ff01011300008067010101130081240300c120830000001300e7a02300176713",
        INIT_15 => X"00276713810007b70007a703810007b702c000ef010104130081242300112623",
        INIT_16 => X"00812623ff01011300008067010101130081240300c120830000001300e7a023",
        INIT_17 => X"00c124030000001300e7a023ff877713810007b70007a703810007b701010413",
        INIT_18 => X"0047f793fec42783fea426230201041300812e23fe0101130000806701010113",
        INIT_19 => X"000080670201011301c124030000001300e7a023fff00713800007b700078863",
        INIT_1A => X"fe040723fcd42823fcc42a23fcb42c23fca42e230301041302812623fd010113",
        INIT_1B => X"fef4478300f70733fdc4270300379793fee447830880006ffe0407a31440006f",
        INIT_1C => X"fef4478300f70733fd84270300379793fee4478300e78023fff0071300f707b3",
        INIT_1D => X"00f707b3fef4478300f70733fd44270300379793fee447830007802300f707b3",
        INIT_1E => X"fff0071300f707b3fef4478300f70733fd04270300379793fee4478300078023",
        INIT_1F => X"00400793f6e7fae300300793fef44703fef407a300178793fef4478300e78023",
        INIT_20 => X"00f707b3fef4478300f70733fdc4270300379793fee447830880006ffef407a3",
        INIT_21 => X"fff0071300f707b3fef4478300f70733fd84270300379793fee4478300078023",
        INIT_22 => X"0007802300f707b3fef4478300f70733fd44270300379793fee4478300e78023",
        INIT_23 => X"00e78023fff0071300f707b3fef4478300f70733fd04270300379793fee44783",
        INIT_24 => X"00178793fee44783f6e7fae300700793fef44703fef407a300178793fef44783",
        INIT_25 => X"fe0407a314c0006ffef4072300400793eae7fce300300793fee44703fef40723",
        INIT_26 => X"0007802300f707b3fef4478300f70733fdc4270300379793fee447830880006f",
        INIT_27 => X"fee447830007802300f707b3fef4478300f70733fd84270300379793fee44783",
        INIT_28 => X"fee4478300e78023fff0071300f707b3fef4478300f70733fd44270300379793",
        INIT_29 => X"fef4478300e78023fff0071300f707b3fef4478300f70733fd04270300379793",
        INIT_2A => X"0900006ffef407a300400793f6e7fae300300793fef44703fef407a300178793",
        INIT_2B => X"00e7802307f0071300f707b3fef4478300f70733fdc4270300379793fee44783",
        INIT_2C => X"00e7802307f0071300f707b3fef4478300f70733fd84270300379793fee44783",
        INIT_2D => X"00e7802307f0071300f707b3fef4478300f70733fd44270300379793fee44783",
        INIT_2E => X"00e78023fff0071300f707b3fef4478300f70733fd04270300379793fee44783",
        INIT_2F => X"00178793fee44783f6e7f6e300700793fef44703fef407a300178793fef44783",
        INIT_30 => X"0301011302c124030000001300000013eae7f8e300700793fee44703fef40723",
        INIT_31 => X"0380006ffe042623fcb42c23fca42e230301041302812623fd01011300008067",
        INIT_32 => X"fdc42783fef4262300f707b3fdc42783fec4270300078a630017f793fd842783",
        INIT_33 => X"fec42783fc0794e3fd842783fcf42c230017d793fd842783fcf42e2300179793",
        INIT_34 => X"fca42c230301041302812623fd010113000080670301011302c1240300078513",
        INIT_35 => X"fd84260301869693fdc42683fed407a300168693fef44683fe0407a3fcb42e23",
        INIT_36 => X"fdc42603fd842683fcf42e23fce42c230086d793fdc4268300e6e73300865713",
        INIT_37 => X"fd010113000080670301011302c1240300078513fef44783fc0692e300c6e6b3",
        INIT_38 => X"00369693fd744683fcd40ba300060693fcb42e23fca42c230301041302812623",
        INIT_39 => X"0006ca63fe068693fec426830d00006ffed42623ff868693fe842683fed42423",
        INIT_3A => X"fec4268301f0059300169613fdc426830380006f0000079300d65733fdc42603",
        INIT_3B => X"fdc42603fec4268300e6e73300c5d733fd842583fec4260300d616b340d586b3",
        INIT_3C => X"000685934106c683000026b7fed422230ff6f693fe442683fee4222300d657b3",
        INIT_3D => X"4106c683000026b700c6802300b686b301068693000026b70ff6f613fe442683",
        INIT_3E => X"000026b700c6a023800006b70006c60300c686b301068693000026b700068613",
        INIT_3F => X"fed42623ff868693fec4268340c68823000026b70ff6f613001686934106c683",
        INIT_40 => X"fe010113000080670301011302c124030000001300000013f206d8e3fec42683",
        INIT_41 => X"00058793fef407a300068713000507930201041300912a2300812c2300112e23",
        INIT_42 => X"0007851300300593fef44783fef4062300070793fef406a300060793fef40723",
        INIT_43 => X"00f484b300050793db1ff0ef0007851300500593fee4478300050493dc5ff0ef",
        INIT_44 => X"00b00593fec4478300f484b300050793d99ff0ef0007851300700593fed44783",
        INIT_45 => X"0181240301c120830007851303f7f79300f487b300050793d81ff0ef00078513",
        INIT_46 => X"00058713000507930301041302812623fd010113000080670201011301412483",
        INIT_47 => X"0ff7f79340f707b3fde4478300078713fdf44783fcf40f2300070793fcf40fa3",
        INIT_48 => X"00812e23fe010113000080670301011302c1240300078513fef44783fef407a3",
        INIT_49 => X"0007c70300f707b3fec4278301078713000027b702c0006ffe04262302010413",
        INIT_4A => X"000787134107c783000027b7fef4262300178793fec4278300e7a023800007b7",
        INIT_4B => X"d4010113000080670201011301c124030000001300000013fce7c4e3fec42783",
        INIT_4C => X"2b7120232b6122232b5124232b4126232b3128232b212a232a812c232a112e23",
        INIT_4D => X"fc0406a3fc040723fc0407a32c01041329b1282329a12a2329912c2329812e23",
        INIT_4E => X"ee840713ea840613e6840693fc042023fcf405a3fff00793fcf40623fff00793",
        INIT_4F => X"00279793fbc427830240006ffa042e23955ff0ef0007851300070593f2840793",
        INIT_50 => X"03f00793fbc42703faf42e2300178793fbc42783d807ac23008787b3fd078793",
        INIT_51 => X"00078713000027b7000786934107c783000027b707c0006ffa042c23fce7dce3",
        INIT_52 => X"000027b700e7802300d787b301078793000027b70007c70300f707b3fb842783",
        INIT_53 => X"00e7a023800007b70007c70300e787b301078793000027b7000787134107c783",
        INIT_54 => X"00178793fb84278340e78823000027b70ff7f713001787934107c783000027b7",
        INIT_55 => X"d4f42c230047a78300078793000027b7f8e7d0e300300793fb842703faf42c23",
        INIT_56 => X"0087a78300078793000027b7c2dff0efd5c42583d584250300400613d4042e23",
        INIT_57 => X"00078793000027b7c09ff0efd5442583d504250300400613d4042a23d4f42823",
        INIT_58 => X"000027b7be5ff0efd4c42583d484250300100613d4042623d4f4242300c7c783",
        INIT_59 => X"bc1ff0ef000d8593000d05130010061300000d9300078d1300d7c78300078793",
        INIT_5A => X"0040079300c7c70300078793000027b75d00006ffa040b235f00006ffa040ba3",
        INIT_5B => X"f587c78300e787b3008787b3fd07879300379793fb644703fb74478308f71a63",
        INIT_5C => X"f187c78300d787b3008787b3fd07879300379793fb644683fb74478301879713",
        INIT_5D => X"00d787b3008787b3fd07879300379793fb644683fb74478300f7673301079793",
        INIT_5E => X"008787b3fd07879300379793fb644683fb74478300f7673300879793ed87c783",
        INIT_5F => X"00379793fb644703fb74478306c0006ffcf4222300f767b3e987c78300d787b3",
        INIT_60 => X"00379793fb644683fb74478301079713f587c78300e787b3008787b3fd078793",
        INIT_61 => X"fb644683fb74478300f7673300879793f187c78300d787b3008787b3fd078793",
        INIT_62 => X"fc442703fcf4222300f767b3ed87c78300d787b3008787b3fd07879300379793",
        INIT_63 => X"40c0006ffcf405a30ff7f793001787930ff7f793fcb4078300f71e63fc042783",
        INIT_64 => X"f8f42c230c078793fcb4078304f7106303e00793fcb407030007d863fcb40783",
        INIT_65 => X"f984250300078613000507939e1ff0eff9c42583f9842503f8f42e2341f7d793",
        INIT_66 => X"fd07879300379793fb644703fb744783fcf405a3fff00793a39ff0eff9c42583",
        INIT_67 => X"008787b3fd07879300379793fb644703fb744783f587c50300e787b3008787b3",
        INIT_68 => X"00e787b3008787b3fd07879300379793fb644703fb744783f187c58300e787b3",
        INIT_69 => X"e987c78300e787b3008787b3fd07879300379793fb644703fb744783ed87c603",
        INIT_6A => X"008787b3fd07879300279793f9744783f8f40ba300050793ad9ff0ef00078693",
        INIT_6B => X"f6842503f6042623f6f424230ff7f793f974478302f71c63fc442703d987a783",
        INIT_6C => X"2ec0006f965ff0eff6c42583f6842503000786130005079390dff0eff6c42583",
        INIT_6D => X"fb644703fb744783d8e7ac23fc442703008787b3fd07879300279793f9744783",
        INIT_6E => X"0007851300070593fcf44703f587c78300e787b3008787b3fd07879300379793",
        INIT_6F => X"008787b3fd07879300379793fb644703fb744783f8f40b2300050793aedff0ef",
        INIT_70 => X"f8f40aa300050793ab9ff0ef0007851300070593fce44703f187c78300e787b3",
        INIT_71 => X"fcd44703ed87c78300e787b3008787b3fd07879300379793fb644703fb744783",
        INIT_72 => X"0cf74063ffe00793f9640703f8f40a2300050793a85ff0ef0007851300070593",
        INIT_73 => X"00100793f95407030af74463ffe00793f95407030ae7ca6300100793f9640703",
        INIT_74 => X"fb74478308e7c26300100793f944070308f74863ffe00793f944070308e7ce63",
        INIT_75 => X"06f71063fcc44703e987c78300e787b3008787b3fd07879300379793fb644703",
        INIT_76 => X"00f767330027979300278793f95407830407e7130047979300278793f9640783",
        INIT_77 => X"f8c42583f8842503f8f4262341f7d793f8f4242300f767b300278793f9440783",
        INIT_78 => X"f95407031700006ffe8ff0eff8c42583f88425030007861300050793f90ff0ef",
        INIT_79 => X"40f70733f9540783f96407030ee7c46301f00793f95407030ef74a63fe000793",
        INIT_7A => X"f94407030ce7c0630070079340f70733f9540783f96407030cf74a63ff800793",
        INIT_7B => X"0040079340f70733f9540783f94407030af74663ffc0079340f70733f9540783",
        INIT_7C => X"e987c78300e787b3008787b3fd07879300379793fb644703fb74478308e7cc63",
        INIT_7D => X"f964068300f76733000087b70087971302078793f954078306f71a63fcc44703",
        INIT_7E => X"40f687b3f9540783f944068300f76733004797930087879340f687b3f9540783",
        INIT_7F => X"e94ff0eff8442583f8042503f8f4222341f7d793f8f4202300f767b300878793",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"00078793000027b70740006feecff0eff8442583f80425030007861300050793",
        INIT_01 => X"0ff9eb9300096b130000099300078913fc44278302f71a630040079300c7c703",
        INIT_02 => X"fc4427830300006fea8ff0eff7442583f704250300500613f7742a23f7642823",
        INIT_03 => X"f784250300400613f7942e23f7842c230feaec93000a6c1300000a9300078a13",
        INIT_04 => X"fd07879300379793fb644703fb744783fcf42023fc442783e78ff0eff7c42583",
        INIT_05 => X"fd07879300379793fb644703fb744783fcf407a3f587c78300e787b3008787b3",
        INIT_06 => X"fd07879300379793fb644703fb744783fcf40723f187c78300e787b3008787b3",
        INIT_07 => X"fd07879300379793fb644703fb744783fcf406a3ed87c78300e787b3008787b3",
        INIT_08 => X"fb644703faf40b2300178793fb644783fcf40623e987c78300e787b3008787b3",
        INIT_09 => X"a0e7f6e300700793fb744703faf40ba300178793fb744783a2e7f6e300700793",
        INIT_0A => X"faf424230c078793fcb4078304f7106303e00793fcb407030007d863fcb40783",
        INIT_0B => X"fa8425030007861300050793d20ff0effac42583fa842503faf4262341f7d793",
        INIT_0C => X"faf42223fae420230000079300100713fcf405a3fff00793d78ff0effac42583",
        INIT_0D => X"2b8124032bc120830007851300000793d50ff0effa442583fa04250300800613",
        INIT_0E => X"29812c8329c12c032a012b832a412b032a812a832ac12a032b0129832b412903",
        INIT_0F => X"00000000000000000000000000000000000080672c01011329012d8329412d03",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;

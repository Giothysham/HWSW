--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"005126230041242300312223001120230000001300000013000000131080006f",
        INIT_01 => X"02d1262302c1242302b1222302a1202300912e2300812c2300712a2300612823",
        INIT_02 => X"0551262305412423053122230521202303112e2303012c2302f12a2302e12823",
        INIT_03 => X"07d1262307c1242307b1222307a1202305912e2305812c2305712a2305612823",
        INIT_04 => X"0101230300c12283008122030041218300012083270000ef07f12a2307e12823",
        INIT_05 => X"0301270302c1268302812603024125830201250301c124830181240301412383",
        INIT_06 => X"05012b0304c12a8304812a03044129830401290303c128830381280303412783",
        INIT_07 => X"07012f0306c12e8306812e0306412d8306012d0305c12c8305812c0305412b83",
        INIT_08 => X"0000031300000293000002130000019300000113000000933020007307412f83",
        INIT_09 => X"0000071300000693000006130000059300000513000004930000041300000393",
        INIT_0A => X"00000b1300000a9300000a130000099300000913000008930000081300000793",
        INIT_0B => X"00000f1300000e9300000e1300000d9300000d1300000c9300000c1300000b93",
        INIT_0C => X"000101130000113700018213eef18193deadc1b7fe0101130000113700000f93",
        INIT_0D => X"ff4101130540006f794000ef0010007379c000effff00113e701011300000117",
        INIT_0E => X"00029663fff50293000583330280006f00051463006124230051222300112023",
        INIT_0F => X"004122830001208300030533fe029ce3fff2829300b303330140006f00058533",
        INIT_10 => X"0000000000000000000000000000006f0000006f0000806700c1011300812303",
        INIT_11 => X"00e7a02300776713810007b70007a703810007b70101041300812623ff010113",
        INIT_12 => X"010104130081242300112623ff010113000080670101011300c1240300000013",
        INIT_13 => X"00c120830000001300e7a02300176713810007b70007a703810007b7068000ef",
        INIT_14 => X"02c000ef010104130081242300112623ff010113000080670101011300812403",
        INIT_15 => X"0081240300c120830000001300e7a02300276713810007b70007a703810007b7",
        INIT_16 => X"810007b70007a703810007b70101041300812623ff0101130000806701010113",
        INIT_17 => X"00812e23fe010113000080670101011300c124030000001300e7a023ff877713",
        INIT_18 => X"00e7a023fff00713800007b7000788630047f793fec42783fea4262302010413",
        INIT_19 => X"fca42e230301041302812623fd010113000080670201011301c1240300000013",
        INIT_1A => X"fee447830880006ffe0407a31440006ffe040723fcd42823fcc42a23fcb42c23",
        INIT_1B => X"fee4478300e78023fff0071300f707b3fef4478300f70733fdc4270300379793",
        INIT_1C => X"00379793fee447830007802300f707b3fef4478300f70733fd84270300379793",
        INIT_1D => X"fd04270300379793fee447830007802300f707b3fef4478300f70733fd442703",
        INIT_1E => X"fef407a300178793fef4478300e78023fff0071300f707b3fef4478300f70733",
        INIT_1F => X"00379793fee447830880006ffef407a300400793f6e7fae300300793fef44703",
        INIT_20 => X"fd84270300379793fee447830007802300f707b3fef4478300f70733fdc42703",
        INIT_21 => X"fd44270300379793fee4478300e78023fff0071300f707b3fef4478300f70733",
        INIT_22 => X"00f70733fd04270300379793fee447830007802300f707b3fef4478300f70733",
        INIT_23 => X"fef44703fef407a300178793fef4478300e78023fff0071300f707b3fef44783",
        INIT_24 => X"eae7fce300300793fee44703fef4072300178793fee44783f6e7fae300700793",
        INIT_25 => X"fdc4270300379793fee447830880006ffe0407a314c0006ffef4072300400793",
        INIT_26 => X"00f70733fd84270300379793fee447830007802300f707b3fef4478300f70733",
        INIT_27 => X"fef4478300f70733fd44270300379793fee447830007802300f707b3fef44783",
        INIT_28 => X"fef4478300f70733fd04270300379793fee4478300e78023fff0071300f707b3",
        INIT_29 => X"00300793fef44703fef407a300178793fef4478300e78023fff0071300f707b3",
        INIT_2A => X"00f70733fdc4270300379793fee447830900006ffef407a300400793f6e7fae3",
        INIT_2B => X"00f70733fd84270300379793fee4478300e7802307f0071300f707b3fef44783",
        INIT_2C => X"00f70733fd44270300379793fee4478300e7802307f0071300f707b3fef44783",
        INIT_2D => X"00f70733fd04270300379793fee4478300e7802307f0071300f707b3fef44783",
        INIT_2E => X"fef44703fef407a300178793fef4478300e78023fff0071300f707b3fef44783",
        INIT_2F => X"eae7f8e300700793fee44703fef4072300178793fee44783f6e7f6e300700793",
        INIT_30 => X"0301041302812623fd010113000080670301011302c124030000001300000013",
        INIT_31 => X"fec4270300078a630017f793fd8427830380006ffe042623fcb42c23fca42e23",
        INIT_32 => X"0017d793fd842783fcf42e2300179793fdc42783fef4262300f707b3fdc42783",
        INIT_33 => X"000080670301011302c1240300078513fec42783fc0794e3fd842783fcf42c23",
        INIT_34 => X"00168693fef44683fe0407a3fcb42e23fca42c230301041302812623fd010113",
        INIT_35 => X"0086d793fdc4268300e6e73300865713fd84260301869693fdc42683fed407a3",
        INIT_36 => X"00078513fef44783fc0692e300c6e6b3fdc42603fd842683fcf42e23fce42c23",
        INIT_37 => X"fcb42e23fca42c230301041302812623fd010113000080670301011302c12403",
        INIT_38 => X"fed42623ff868693fe842683fed4242300369693fd744683fcd40ba300060693",
        INIT_39 => X"0380006f0000079300d65733fdc426030006ca63fe068693fec426830ac0006f",
        INIT_3A => X"fd842583fec4260300d616b340d586b3fec4268301f0059300169613fdc42683",
        INIT_3B => X"0ff6f693fe442683fee4222300d657b3fdc42603fec4268300e6e73300c5d733",
        INIT_3C => X"01068693000026b70ff6f613fe442683000685934106c683000026b7fed42223",
        INIT_3D => X"40c68823000026b70ff6f613001686934106c683000026b700c6802300b686b3",
        INIT_3E => X"02c124030000001300000013f406dae3fec42683fed42623ff868693fec42683",
        INIT_3F => X"000507930201041300912a2300812c2300112e23fe0101130000806703010113",
        INIT_40 => X"fef4062300070793fef406a300060793fef4072300058793fef407a300068713",
        INIT_41 => X"0007851300500593fee4478300050493de9ff0ef0007851300300593fef44783",
        INIT_42 => X"00050793dbdff0ef0007851300700593fed4478300f484b300050793dd5ff0ef",
        INIT_43 => X"03f7f79300f487b300050793da5ff0ef0007851300b00593fec4478300f484b3",
        INIT_44 => X"02812623fd0101130000806702010113014124830181240301c1208300078513",
        INIT_45 => X"00078713fdf44783fcf40f2300070793fcf40fa3000587130005079303010413",
        INIT_46 => X"0301011302c1240300078513fef44783fef407a30ff7f79340f707b3fde44783",
        INIT_47 => X"01078713000027b702c0006ffe0426230201041300812e23fe01011300008067",
        INIT_48 => X"fef4262300178793fec4278300e7a023800007b70007c70300f707b3fec42783",
        INIT_49 => X"01c124030000001300000013fce7c4e3fec42783000787134107c783000027b7",
        INIT_4A => X"2b4126232b3128232b212a232a812c232a112e23d40101130000806702010113",
        INIT_4B => X"2c01041329b1282329a12a2329912c2329812e232b7120232b6122232b512423",
        INIT_4C => X"fc042023fcf405a3fff00793fcf40623fff00793fc0406a3fc040723fc0407a3",
        INIT_4D => X"fa042e23979ff0ef0007851300070593f2840793ee840713ea840613e6840693",
        INIT_4E => X"00178793fbc42783d807ac23008787b3fd07879300279793fbc427830240006f",
        INIT_4F => X"4107c783000027b70580006ffa042c23fce7dce303f00793fbc42703faf42e23",
        INIT_50 => X"01078793000027b70007c70300f707b3fb84278300078713000027b700078693",
        INIT_51 => X"40e78823000027b70ff7f713001787934107c783000027b700e7802300d787b3",
        INIT_52 => X"00078793000027b7fae7d2e300300793fb842703faf42c2300178793fb842783",
        INIT_53 => X"000027b7c75ff0efd5c42583d584250300400613d4042e23d4f42c230047a783",
        INIT_54 => X"c51ff0efd5442583d504250300400613d4042a23d4f428230087a78300078793",
        INIT_55 => X"d4c42583d484250300100613d4042623d4f4242300c7c78300078793000027b7",
        INIT_56 => X"000d05130010061300000d9300078d1300d7c78300078793000027b7c2dff0ef",
        INIT_57 => X"00078793000027b75d00006ffa040b235f00006ffa040ba3c09ff0ef000d8593",
        INIT_58 => X"008787b3fd07879300379793fb644703fb74478308f71a630040079300c7c703",
        INIT_59 => X"008787b3fd07879300379793fb644683fb74478301879713f587c78300e787b3",
        INIT_5A => X"fd07879300379793fb644683fb74478300f7673301079793f187c78300d787b3",
        INIT_5B => X"00379793fb644683fb74478300f7673300879793ed87c78300d787b3008787b3",
        INIT_5C => X"fb74478306c0006ffcf4222300f767b3e987c78300d787b3008787b3fd078793",
        INIT_5D => X"fb74478301079713f587c78300e787b3008787b3fd07879300379793fb644703",
        INIT_5E => X"00f7673300879793f187c78300d787b3008787b3fd07879300379793fb644683",
        INIT_5F => X"00f767b3ed87c78300d787b3008787b3fd07879300379793fb644683fb744783",
        INIT_60 => X"0ff7f793001787930ff7f793fcb4078300f71e63fc042783fc442703fcf42223",
        INIT_61 => X"fcb4078304f7106303e00793fcb407030007d863fcb4078340c0006ffcf405a3",
        INIT_62 => X"00050793a29ff0eff9c42583f9842503f8f42e2341f7d793f8f42c230c078793",
        INIT_63 => X"fb644703fb744783fcf405a3fff00793a81ff0eff9c42583f984250300078613",
        INIT_64 => X"00379793fb644703fb744783f587c50300e787b3008787b3fd07879300379793",
        INIT_65 => X"fd07879300379793fb644703fb744783f187c58300e787b3008787b3fd078793",
        INIT_66 => X"008787b3fd07879300379793fb644703fb744783ed87c60300e787b3008787b3",
        INIT_67 => X"00279793f9744783f8f40ba300050793afdff0ef00078693e987c78300e787b3",
        INIT_68 => X"f6f424230ff7f793f974478302f71c63fc442703d987a783008787b3fd078793",
        INIT_69 => X"f6c42583f68425030007861300050793955ff0eff6c42583f6842503f6042623",
        INIT_6A => X"d8e7ac23fc442703008787b3fd07879300279793f97447832ec0006f9adff0ef",
        INIT_6B => X"fcf44703f587c78300e787b3008787b3fd07879300379793fb644703fb744783",
        INIT_6C => X"00379793fb644703fb744783f8f40b2300050793b11ff0ef0007851300070593",
        INIT_6D => X"addff0ef0007851300070593fce44703f187c78300e787b3008787b3fd078793",
        INIT_6E => X"00e787b3008787b3fd07879300379793fb644703fb744783f8f40aa300050793",
        INIT_6F => X"f9640703f8f40a2300050793aa9ff0ef0007851300070593fcd44703ed87c783",
        INIT_70 => X"0af74463ffe00793f95407030ae7ca6300100793f96407030cf74063ffe00793",
        INIT_71 => X"00100793f944070308f74863ffe00793f944070308e7ce6300100793f9540703",
        INIT_72 => X"e987c78300e787b3008787b3fd07879300379793fb644703fb74478308e7c263",
        INIT_73 => X"00278793f95407830407e7130047979300278793f964078306f71063fcc44703",
        INIT_74 => X"f8f4262341f7d793f8f4242300f767b300278793f944078300f7673300279793",
        INIT_75 => X"831ff0eff8c42583f88425030007861300050793fd8ff0eff8c42583f8842503",
        INIT_76 => X"f96407030ee7c46301f00793f95407030ef74a63fe000793f95407031700006f",
        INIT_77 => X"0070079340f70733f9540783f96407030cf74a63ff80079340f70733f9540783",
        INIT_78 => X"f9540783f94407030af74663ffc0079340f70733f9540783f94407030ce7c063",
        INIT_79 => X"008787b3fd07879300379793fb644703fb74478308e7cc630040079340f70733",
        INIT_7A => X"000087b70087971302078793f954078306f71a63fcc44703e987c78300e787b3",
        INIT_7B => X"f944068300f76733004797930087879340f687b3f9540783f964068300f76733",
        INIT_7C => X"f8042503f8f4222341f7d793f8f4202300f767b30087879340f687b3f9540783",
        INIT_7D => X"0740006ff34ff0eff8442583f80425030007861300050793edcff0eff8442583",
        INIT_7E => X"0000099300078913fc44278302f71a630040079300c7c70300078793000027b7",
        INIT_7F => X"ef0ff0eff7442583f704250300500613f7742a23f76428230ff9eb9300096b13",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"f7942e23f7842c230feaec93000a6c1300000a9300078a13fc4427830300006f",
        INIT_01 => X"fb644703fb744783fcf42023fc442783ec0ff0eff7c42583f784250300400613",
        INIT_02 => X"fb644703fb744783fcf407a3f587c78300e787b3008787b3fd07879300379793",
        INIT_03 => X"fb644703fb744783fcf40723f187c78300e787b3008787b3fd07879300379793",
        INIT_04 => X"fb644703fb744783fcf406a3ed87c78300e787b3008787b3fd07879300379793",
        INIT_05 => X"00178793fb644783fcf40623e987c78300e787b3008787b3fd07879300379793",
        INIT_06 => X"fb744703faf40ba300178793fb744783a2e7f6e300700793fb644703faf40b23",
        INIT_07 => X"fcb4078304f7106303e00793fcb407030007d863fcb40783a0e7f6e300700793",
        INIT_08 => X"00050793d68ff0effac42583fa842503faf4262341f7d793faf424230c078793",
        INIT_09 => X"0000079300100713fcf405a3fff00793dc0ff0effac42583fa84250300078613",
        INIT_0A => X"00000793f8cff0efd98ff0effa442583fa04250300800613faf42223fae42023",
        INIT_0B => X"2a412b032a812a832ac12a032b0129832b4129032b8124032bc1208300078513",
        INIT_0C => X"00000000000080672c01011329012d8329412d0329812c8329c12c032a012b83",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;

--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"0000041300000393000003130000029300000213000001930000011300000093",
        INIT_01 => X"0000081300000793000007130000069300000613000005930000051300000493",
        INIT_02 => X"00000c1300000b9300000b1300000a9300000a13000009930000091300000893",
        INIT_03 => X"0000113700000f9300000f1300000e9300000e1300000d9300000d1300000c93",
        INIT_04 => X"3004507334011073000101130000113700018213eef18193deadc1b7fe010113",
        INIT_05 => X"00112023ff4101130540006f6fc000ef00100073704000ef30411073fff00113",
        INIT_06 => X"0005853300029663fff50293000583330280006f000514630061242300512223",
        INIT_07 => X"00812303004122830001208300030533fe029ce3fff2829300b303330140006f",
        INIT_08 => X"810007b70101041300812623ff0101130000006f0000006f0000806700c10113",
        INIT_09 => X"000080670101011300c124030000001300e7a02300776713810007b70007a703",
        INIT_0A => X"810007b70007a703810007b7068000ef010104130081242300112623ff010113",
        INIT_0B => X"ff01011300008067010101130081240300c120830000001300e7a02300176713",
        INIT_0C => X"00276713810007b70007a703810007b702c000ef010104130081242300112623",
        INIT_0D => X"00812623ff01011300008067010101130081240300c120830000001300e7a023",
        INIT_0E => X"00c124030000001300e7a023ff877713810007b70007a703810007b701010413",
        INIT_0F => X"00100713000027b7fea426230201041300812e23fe0101130000806701010113",
        INIT_10 => X"0000001300e7a02300700713810007b700e7a02301700713810007b700e7aa23",
        INIT_11 => X"fcb42c23fca42e230301041302812623fd010113000080670201011301c12403",
        INIT_12 => X"00179793fee447830880006ffe0407a31400006ffe040723fcd42823fcc42a23",
        INIT_13 => X"00179793fee4478300e78023fff0071300f707b3fef4478300f70733fdc42703",
        INIT_14 => X"fd44270300179793fee447830007802300f707b3fef4478300f70733fd842703",
        INIT_15 => X"00f70733fd04270300179793fee447830007802300f707b3fef4478300f70733",
        INIT_16 => X"fef44783fef407a300178793fef4478300e78023fff0071300f707b3fef44783",
        INIT_17 => X"00f70733fdc4270300179793fee447830880006ffef407a300100793f6078ce3",
        INIT_18 => X"fef4478300f70733fd84270300179793fee447830007802300f707b3fef44783",
        INIT_19 => X"fef4478300f70733fd44270300179793fee4478300e78023fff0071300f707b3",
        INIT_1A => X"00f707b3fef4478300f70733fd04270300179793fee447830007802300f707b3",
        INIT_1B => X"f6e7fae300100793fef44703fef407a300178793fef4478300e78023fff00713",
        INIT_1C => X"1480006ffef4072300100793ec0780e3fee44783fef4072300178793fee44783",
        INIT_1D => X"00f707b3fef4478300f70733fdc4270300179793fee447830880006ffe0407a3",
        INIT_1E => X"0007802300f707b3fef4478300f70733fd84270300179793fee4478300078023",
        INIT_1F => X"00e78023fff0071300f707b3fef4478300f70733fd44270300179793fee44783",
        INIT_20 => X"00e78023fff0071300f707b3fef4478300f70733fd04270300179793fee44783",
        INIT_21 => X"0900006ffef407a300100793f6078ce3fef44783fef407a300178793fef44783",
        INIT_22 => X"00e7802307f0071300f707b3fef4478300f70733fdc4270300179793fee44783",
        INIT_23 => X"00e7802307f0071300f707b3fef4478300f70733fd84270300179793fee44783",
        INIT_24 => X"00e7802307f0071300f707b3fef4478300f70733fd44270300179793fee44783",
        INIT_25 => X"00e78023fff0071300f707b3fef4478300f70733fd04270300179793fee44783",
        INIT_26 => X"00178793fee44783f6e7f6e300100793fef44703fef407a300178793fef44783",
        INIT_27 => X"0301011302c124030000001300000013eae7fae300100793fee44703fef40723",
        INIT_28 => X"0380006ffe042623fcb42c23fca42e230301041302812623fd01011300008067",
        INIT_29 => X"fdc42783fef4262300f707b3fdc42783fec4270300078a630017f793fd842783",
        INIT_2A => X"fec42783fc0794e3fd842783fcf42c230017d793fd842783fcf42e2300179793",
        INIT_2B => X"fca42e230301041302812623fd010113000080670301011302c1240300078513",
        INIT_2C => X"fdc42783fcf42e234087d793fdc42783fef4262300178793fec42783fe042623",
        INIT_2D => X"02812623fd010113000080670301011302c1240300078513fec42783fe0792e3",
        INIT_2E => X"fe842683fed4242300369693fd442683fcc42a23fcb42e23fca42c2303010413",
        INIT_2F => X"00d65733fdc426030006ca63fe068693fec426830ac0006ffed42623ff868693",
        INIT_30 => X"00d616b340d586b3fec4268301f0059300169613fdc426830380006f00000793",
        INIT_31 => X"fee4222300d657b3fdc42603fec4268300e6e73300c5d733fd842583fec42603",
        INIT_32 => X"00d606b3800006b7000686130106c683000026b7fed422230ff6f693fe442683",
        INIT_33 => X"0ff6f613001686930106c683000026b700d600230ff6f693fe44268300068613",
        INIT_34 => X"00000013f406dae3fec42683fed42623ff868693fec4268300c68823000026b7",
        INIT_35 => X"00912a2300812c2300112e23fe010113000080670301011302c1240300000013",
        INIT_36 => X"fef406a300060793fef4072300058793fef407a3000687130005079302010413",
        INIT_37 => X"fee4478300050493e11ff0ef0007851300300593fef44783fef4062300070793",
        INIT_38 => X"0007851300700593fed4478300f484b300050793dfdff0ef0007851300500593",
        INIT_39 => X"00050793dcdff0ef0007851300b00593fec4478300f484b300050793de5ff0ef",
        INIT_3A => X"0000806702010113014124830181240301c120830007851303f7f79300f487b3",
        INIT_3B => X"fcf40f2300070793fcf40fa300058713000507930301041302812623fd010113",
        INIT_3C => X"00078513fef44783fef407a30ff7f79340f707b3fde4478300078713fdf44783",
        INIT_3D => X"1b3128231b212a231a812c231a112e23e4010113000080670301011302c12403",
        INIT_3E => X"19b1282319a12a2319912c2319812e231b7120231b6122231b5124231b412623",
        INIT_3F => X"fcf405a3fff00793fcf40623fff00793fc0406a3fc040723fc0407a31c010413",
        INIT_40 => X"a11ff0ef0007851300070593f6c40793f6840713f6440613f6040693fc042023",
        INIT_41 => X"fbf44783e807a823008787b3fd07879300279793fbf447830240006ffa040fa3",
        INIT_42 => X"fbe447830580006ffa040f23fce7fce303f00793fbf44703faf40fa300178793",
        INIT_43 => X"00070713000027370007069300e6873380000737000706930107470300002737",
        INIT_44 => X"000027b70ff7f713001787930107c783000027b700f680230007c78300f707b3",
        INIT_45 => X"000027b7fae7f2e300300793fbe44703faf40f2300178793fbe4478300e78823",
        INIT_46 => X"cddff0efe5c42583e584250300400613e4042e23e4f42c230047a78300078793",
        INIT_47 => X"e5442583e504250300400613e4042a23e4f428230087a78300078793000027b7",
        INIT_48 => X"e484250300100613e4042623e4f4242300c7c78300078793000027b7cb9ff0ef",
        INIT_49 => X"0010061300000d9300078d1300d7c78300078793000027b7c95ff0efe4c42583",
        INIT_4A => X"000027b75d00006ffa040e235f00006ffa040ea3c71ff0ef000d8593000d0513",
        INIT_4B => X"fd07879300179793fbc44703fbd4478308f71a630040079300c7c70300078793",
        INIT_4C => X"fd07879300179793fbc44683fbd4478301879713f9c7c78300e787b3008787b3",
        INIT_4D => X"00179793fbc44683fbd4478300f7673301079793f987c78300d787b3008787b3",
        INIT_4E => X"fbc44683fbd4478300f7673300879793f947c78300d787b3008787b3fd078793",
        INIT_4F => X"06c0006ffcf4222300f767b3f907c78300d787b3008787b3fd07879300179793",
        INIT_50 => X"01079713f9c7c78300e787b3008787b3fd07879300179793fbc44703fbd44783",
        INIT_51 => X"00879793f987c78300d787b3008787b3fd07879300179793fbc44683fbd44783",
        INIT_52 => X"f947c78300d787b3008787b3fd07879300179793fbc44683fbd4478300f76733",
        INIT_53 => X"001787930ff7f793fcb4078300f71e63fc042783fc442703fcf4222300f767b3",
        INIT_54 => X"04f7106303e00793fcb407030007d863fcb4078340c0006ffcf405a30ff7f793",
        INIT_55 => X"ab5ff0ef00078513fa042783faf4222341f7d793faf420230c078793fcb40783",
        INIT_56 => X"fbd44783fcf405a3fff00793ae9ff0effa442583fa0425030007861300050793",
        INIT_57 => X"fbc44703fbd44783f9c7c50300e787b3008787b3fd07879300179793fbc44703",
        INIT_58 => X"00179793fbc44703fbd44783f987c58300e787b3008787b3fd07879300179793",
        INIT_59 => X"fd07879300179793fbc44703fbd44783f947c60300e787b3008787b3fd078793",
        INIT_5A => X"f9f44783f8f40fa300050793b61ff0ef00078693f907c78300e787b3008787b3",
        INIT_5B => X"0ff7f793f9f4478302f71c63fc442703e907a783008787b3fd07879300279793",
        INIT_5C => X"f704250300078613000507939e1ff0ef00078513f7042783f6042a23f6f42823",
        INIT_5D => X"fc442703008787b3fd07879300279793f9f447832ec0006fa15ff0eff7442583",
        INIT_5E => X"f9c7c78300e787b3008787b3fd07879300179793fbc44703fbd44783e8e7a823",
        INIT_5F => X"fbc44703fbd44783f8f40f2300050793b75ff0ef0007851300070593fcf44703",
        INIT_60 => X"0007851300070593fce44703f987c78300e787b3008787b3fd07879300179793",
        INIT_61 => X"008787b3fd07879300179793fbc44703fbd44783f8f40ea300050793b41ff0ef",
        INIT_62 => X"f8f40e2300050793b0dff0ef0007851300070593fcd44703f947c78300e787b3",
        INIT_63 => X"ffe00793f9d407030ae7ca6300100793f9e407030cf74063ffe00793f9e40703",
        INIT_64 => X"f9c4070308f74863ffe00793f9c4070308e7ce6300100793f9d407030af74463",
        INIT_65 => X"00e787b3008787b3fd07879300179793fbc44703fbd4478308e7c26300100793",
        INIT_66 => X"f9d407830407e7130047979300278793f9e4078306f71063fcc44703f907c783",
        INIT_67 => X"41f7d793f8f4282300f767b300278793f9c4078300f767330027979300278793",
        INIT_68 => X"f9442583f90425030007861300050793865ff0ef00078513f9042783f8f42a23",
        INIT_69 => X"0ee7c46301f00793f9d407030ef74a63fe000793f9d407031700006f899ff0ef",
        INIT_6A => X"40f70733f9d40783f9e407030cf74a63ff80079340f70733f9d40783f9e40703",
        INIT_6B => X"f9c407030af74663ffc0079340f70733f9d40783f9c407030ce7c06300700793",
        INIT_6C => X"fd07879300179793fbc44703fbd4478308e7cc630040079340f70733f9d40783",
        INIT_6D => X"0087971302078793f9d4078306f71a63fcc44703f907c78300e787b3008787b3",
        INIT_6E => X"00f76733004797930087879340f687b3f9d40783f9e4068300f76733000087b7",
        INIT_6F => X"f8f4262341f7d793f8f4242300f767b30087879340f687b3f9d40783f9c40683",
        INIT_70 => X"f9cff0eff8c42583f88425030007861300050793f68ff0ef00078513f8842783",
        INIT_71 => X"00078913fc44278302f71a630040079300c7c70300078793000027b70740006f",
        INIT_72 => X"f7c42583f784250300500613f7742e23f7642c230ff9eb9300096b1300000993",
        INIT_73 => X"f98420230feaec93000a6c1300000a9300078a13fc4427830300006ff58ff0ef",
        INIT_74 => X"fbd44783fcf42023fc442783f28ff0eff8442583f804250300400613f9942223",
        INIT_75 => X"fbd44783fcf407a3f9c7c78300e787b3008787b3fd07879300179793fbc44703",
        INIT_76 => X"fbd44783fcf40723f987c78300e787b3008787b3fd07879300179793fbc44703",
        INIT_77 => X"fbd44783fcf406a3f947c78300e787b3008787b3fd07879300179793fbc44703",
        INIT_78 => X"fbc44783fcf40623f907c78300e787b3008787b3fd07879300179793fbc44703",
        INIT_79 => X"faf40ea300178793fbd44783a2e7f6e300100793fbc44703faf40e2300178793",
        INIT_7A => X"04f7106303e00793fcb407030007d863fcb40783a0e7f6e300100793fbd44703",
        INIT_7B => X"df4ff0ef00078513fb042783faf42a2341f7d793faf428230c078793fcb40783",
        INIT_7C => X"00100713fcf405a3fff00793e28ff0effb442583fb0425030007861300050793",
        INIT_7D => X"00000793e00ff0effac42583fa84250300800613faf42623fae4242300000793",
        INIT_7E => X"1a412b031a812a831ac12a031b0129831b4129031b8124031bc1208300078513",
        INIT_7F => X"00000000000080671c01011319012d8319412d0319812c8319c12c031a012b83",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;

--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"0000041300000393000003130000029300000213000001930000011300000093",
        INIT_01 => X"0000081300000793000007130000069300000613000005930000051300000493",
        INIT_02 => X"00000c1300000b9300000b1300000a9300000a13000009930000091300000893",
        INIT_03 => X"0000113700000f9300000f1300000e9300000e1300000d9300000d1300000c93",
        INIT_04 => X"3004507334011073000101130000113700018213eef18193deadc1b7fe010113",
        INIT_05 => X"00112023ff4101130540006f6f4000ef001000736fc000ef30411073fff00113",
        INIT_06 => X"0005853300029663fff50293000583330280006f000514630061242300512223",
        INIT_07 => X"00812303004122830001208300030533fe029ce3fff2829300b303330140006f",
        INIT_08 => X"810007b70101041300812623ff0101130000006f0000006f0000806700c10113",
        INIT_09 => X"000080670101011300c124030000001300e7a02300776713810007b70007a703",
        INIT_0A => X"810007b70007a703810007b7068000ef010104130081242300112623ff010113",
        INIT_0B => X"ff01011300008067010101130081240300c120830000001300e7a02300176713",
        INIT_0C => X"00276713810007b70007a703810007b702c000ef010104130081242300112623",
        INIT_0D => X"00812623ff01011300008067010101130081240300c120830000001300e7a023",
        INIT_0E => X"00c124030000001300e7a023ff877713810007b70007a703810007b701010413",
        INIT_0F => X"00100713000027b7fea426230201041300812e23fe0101130000806701010113",
        INIT_10 => X"0000001300e7a02300700713810007b700e7a02301700713810007b700e7aa23",
        INIT_11 => X"fcb42c23fca42e230301041302812623fd010113000080670201011301c12403",
        INIT_12 => X"00179793fee447830880006ffe0407a31400006ffe040723fcd42823fcc42a23",
        INIT_13 => X"00179793fee4478300e78023fff0071300f707b3fef4478300f70733fdc42703",
        INIT_14 => X"fd44270300179793fee447830007802300f707b3fef4478300f70733fd842703",
        INIT_15 => X"00f70733fd04270300179793fee447830007802300f707b3fef4478300f70733",
        INIT_16 => X"fef44783fef407a300178793fef4478300e78023fff0071300f707b3fef44783",
        INIT_17 => X"00f70733fdc4270300179793fee447830880006ffef407a300100793f6078ce3",
        INIT_18 => X"fef4478300f70733fd84270300179793fee447830007802300f707b3fef44783",
        INIT_19 => X"fef4478300f70733fd44270300179793fee4478300e78023fff0071300f707b3",
        INIT_1A => X"00f707b3fef4478300f70733fd04270300179793fee447830007802300f707b3",
        INIT_1B => X"f6e7fae300100793fef44703fef407a300178793fef4478300e78023fff00713",
        INIT_1C => X"1480006ffef4072300100793ec0780e3fee44783fef4072300178793fee44783",
        INIT_1D => X"00f707b3fef4478300f70733fdc4270300179793fee447830880006ffe0407a3",
        INIT_1E => X"0007802300f707b3fef4478300f70733fd84270300179793fee4478300078023",
        INIT_1F => X"00e78023fff0071300f707b3fef4478300f70733fd44270300179793fee44783",
        INIT_20 => X"00e78023fff0071300f707b3fef4478300f70733fd04270300179793fee44783",
        INIT_21 => X"0900006ffef407a300100793f6078ce3fef44783fef407a300178793fef44783",
        INIT_22 => X"00e7802307f0071300f707b3fef4478300f70733fdc4270300179793fee44783",
        INIT_23 => X"00e7802307f0071300f707b3fef4478300f70733fd84270300179793fee44783",
        INIT_24 => X"00e7802307f0071300f707b3fef4478300f70733fd44270300179793fee44783",
        INIT_25 => X"00e78023fff0071300f707b3fef4478300f70733fd04270300179793fee44783",
        INIT_26 => X"00178793fee44783f6e7f6e300100793fef44703fef407a300178793fef44783",
        INIT_27 => X"0301011302c124030000001300000013eae7fae300100793fee44703fef40723",
        INIT_28 => X"0380006ffe042623fcb42c23fca42e230301041302812623fd01011300008067",
        INIT_29 => X"fdc42783fef4262300f707b3fdc42783fec4270300078a630017f793fd842783",
        INIT_2A => X"fec42783fc0794e3fd842783fcf42c230017d793fd842783fcf42e2300179793",
        INIT_2B => X"fca42e230301041302812623fd010113000080670301011302c1240300078513",
        INIT_2C => X"fdc42783fcf42e234087d793fdc42783fef4262300178793fec42783fe042623",
        INIT_2D => X"02812623fd010113000080670301011302c1240300078513fec42783fe0792e3",
        INIT_2E => X"ff868693fe842683fed4242300369693fd842683fcb42c23fca42e2303010413",
        INIT_2F => X"0005c863fe058593fec425830046a6830006a603fdc426830a80006ffed42623",
        INIT_30 => X"00b515b340b805b3fec4258301f008130016951302c0006f0000079300b6d733",
        INIT_31 => X"0ff6f693fe442683fee4222300b6d7b3fec4258300e5e73300a65733fec42503",
        INIT_32 => X"fe4426830006861300d606b3800006b7000686130106c683000026b7fed42223",
        INIT_33 => X"00c68823000026b70ff6f613001686930106c683000026b700d600230ff6f693",
        INIT_34 => X"02c124030000001300000013f406dce3fec42683fed42623ff868693fec42683",
        INIT_35 => X"000507930201041300912a2300812c2300112e23fe0101130000806703010113",
        INIT_36 => X"fef4062300070793fef406a300060793fef4072300058793fef407a300068713",
        INIT_37 => X"0007851300500593fee4478300050493e19ff0ef0007851300300593fef44783",
        INIT_38 => X"00050793dedff0ef0007851300700593fed4478300f484b300050793e05ff0ef",
        INIT_39 => X"03f7f79300f487b300050793dd5ff0ef0007851300b00593fec4478300f484b3",
        INIT_3A => X"02812623fd0101130000806702010113014124830181240301c1208300078513",
        INIT_3B => X"00078713fdf44783fcf40f2300070793fcf40fa3000587130005079303010413",
        INIT_3C => X"0301011302c1240300078513fef44783fef407a30ff7f79340f707b3fde44783",
        INIT_3D => X"1b5124231b4126231b3128231b212a231a812c231a112e23e401011300008067",
        INIT_3E => X"fc0407a31c01041319b1282319a12a2319912c2319812e231b7120231b612223",
        INIT_3F => X"fa840693fc042023fcf405a3fff00793fcf40623fff00793fc0406a3fc040723",
        INIT_40 => X"0240006ffa040fa3a19ff0ef0007851300070593fb440793fb040713fac40613",
        INIT_41 => X"faf40fa300178793fbf44783ec07ac23008787b3fd07879300279793fbf44783",
        INIT_42 => X"0107470300002737fbe447830580006ffa040f23fce7fce303f00793fbf44703",
        INIT_43 => X"0007c78300f707b300070713000027370007069300e687338000073700070693",
        INIT_44 => X"fbe4478300e78823000027b70ff7f713001787930107c783000027b700f68023",
        INIT_45 => X"00478513000027b700400593fae7f2e300300793fbe44703faf40f2300178793",
        INIT_46 => X"00c78513000027b700100593ce9ff0ef00878513000027b700400593cf9ff0ef",
        INIT_47 => X"fa040e236600006ffa040ea3cc9ff0ef00d78513000027b700100593cd9ff0ef",
        INIT_48 => X"fbc44703fbd4478308f71a630040079300c7c70300078793000027b76400006f",
        INIT_49 => X"fbc44683fbd4478301879713fe47c78300e787b3008787b3fd07879300179793",
        INIT_4A => X"fbd4478300f7673301079793fe07c78300d787b3008787b3fd07879300179793",
        INIT_4B => X"00f7673300879793fdc7c78300d787b3008787b3fd07879300179793fbc44683",
        INIT_4C => X"00f767b3fd87c78300d787b3008787b3fd07879300179793fbc44683fbd44783",
        INIT_4D => X"00e787b3008787b3fd07879300179793fbc44703fbd4478306c0006ffcf42223",
        INIT_4E => X"00d787b3008787b3fd07879300179793fbc44683fbd4478301079713fe47c783",
        INIT_4F => X"008787b3fd07879300179793fbc44683fbd4478300f7673300879793fe07c783",
        INIT_50 => X"fcb4078300f71e63fc042783fc442703fcf4222300f767b3fdc7c78300d787b3",
        INIT_51 => X"fcb407030007d863fcb4078347c0006ffcf405a30ff7f793001787930ff7f793",
        INIT_52 => X"e5842783e4f42e2341f7d793e4f42c230c078793fcb4078304f71c6303e00793",
        INIT_53 => X"af5ff0ef0007851300070793e9c42783e9842703e9042e23e8f42c23e5c42803",
        INIT_54 => X"fbd44783fcf405a3fff00793b29ff0ef0007851300070593e984079300050713",
        INIT_55 => X"fbc44703fbd44783fe47c50300e787b3008787b3fd07879300179793fbc44703",
        INIT_56 => X"00179793fbc44703fbd44783fe07c58300e787b3008787b3fd07879300179793",
        INIT_57 => X"fd07879300179793fbc44703fbd44783fdc7c60300e787b3008787b3fd078793",
        INIT_58 => X"fbb44783faf40da300050793b99ff0ef00078693fd87c78300e787b3008787b3",
        INIT_59 => X"0ff7f793fbb4478304f71863fc442703ed87a783008787b3fd07879300279793",
        INIT_5A => X"e9442783e9042703e9042a23e8f42823e5442803e5042783e4042a23e4f42823",
        INIT_5B => X"a3dff0ef0007851300070593e904079300050713a09ff0ef0007851300070793",
        INIT_5C => X"fbd44783ece7ac23fc442703008787b3fd07879300279793fbb4478332c0006f",
        INIT_5D => X"00070593fcf44703fe47c78300e787b3008787b3fd07879300179793fbc44703",
        INIT_5E => X"fd07879300179793fbc44703fbd44783faf40d2300050793b95ff0ef00078513",
        INIT_5F => X"00050793b61ff0ef0007851300070593fce44703fe07c78300e787b3008787b3",
        INIT_60 => X"fdc7c78300e787b3008787b3fd07879300179793fbc44703fbd44783faf40ca3",
        INIT_61 => X"ffe00793fba40703faf40c2300050793b2dff0ef0007851300070593fcd44703",
        INIT_62 => X"fb9407030cf74063ffe00793fb9407030ce7c66300100793fba407030cf74c63",
        INIT_63 => X"08e7ce6300100793fb8407030af74463ffe00793fb8407030ae7ca6300100793",
        INIT_64 => X"fcc44703fd87c78300e787b3008787b3fd07879300179793fbc44703fbd44783",
        INIT_65 => X"0027979300278793fb9407830407e7130047979300278793fba4078306f71c63",
        INIT_66 => X"e4842783e4f4262341f7d793e4f4242300f767b300278793fb84078300f76733",
        INIT_67 => X"875ff0ef0007851300070793e8c42783e8842703e9042623e8f42423e4c42803",
        INIT_68 => X"fe000793fb9407031980006f8a9ff0ef0007851300070593e884079300050713",
        INIT_69 => X"ff80079340f70733fb940783fba4070310e7c06301f00793fb94070310f74663",
        INIT_6A => X"fb940783fb8407030ce7cc630070079340f70733fb940783fba407030ef74663",
        INIT_6B => X"0ae7c8630040079340f70733fb940783fb8407030cf74263ffc0079340f70733",
        INIT_6C => X"fcc44703fd87c78300e787b3008787b3fd07879300179793fbc44703fbd44783",
        INIT_6D => X"fb940783fba4068300f76733000087b70087971302078793fb94078308f71663",
        INIT_6E => X"0087879340f687b3fb940783fb84068300f76733004797930087879340f687b3",
        INIT_6F => X"e9042223e8f42023e4442803e4042783e4f4222341f7d793e4f4202300f767b3",
        INIT_70 => X"00070593e804079300050713f60ff0ef0007851300070793e8442783e8042703",
        INIT_71 => X"02f71e630040079300c7c70300078793000027b70840006ff94ff0ef00078513",
        INIT_72 => X"e6e42c23000b8793000b07130ff9eb9300096b130000099300078913fc442783",
        INIT_73 => X"00078a13fc4427830380006ff48ff0ef0007851300500593e7840793e6f42e23",
        INIT_74 => X"e7040793e6f42a23e6e42823000c8793000c07130feaec93000a6c1300000a93",
        INIT_75 => X"00179793fbc44703fbd44783fcf42023fc442783f10ff0ef0007851300400593",
        INIT_76 => X"00179793fbc44703fbd44783fcf407a3fe47c78300e787b3008787b3fd078793",
        INIT_77 => X"00179793fbc44703fbd44783fcf40723fe07c78300e787b3008787b3fd078793",
        INIT_78 => X"00179793fbc44703fbd44783fcf406a3fdc7c78300e787b3008787b3fd078793",
        INIT_79 => X"faf40e2300178793fbc44783fcf40623fd87c78300e787b3008787b3fd078793",
        INIT_7A => X"00100793fbd44703faf40ea300178793fbd447839ae7fee300100793fbc44703",
        INIT_7B => X"0c078793fcb4078304f7186303e00793fcb407030007d863fcb4078398e7fee3",
        INIT_7C => X"00070793e6c42783e6842703e7b42623e7a4242300078d9341f7d79300078d13",
        INIT_7D => X"fff00793e00ff0ef0007851300070593e684079300050713dccff0ef00078513",
        INIT_7E => X"0007851300800593ea040793eaf42223eae420230000079300100713fcf405a3",
        INIT_7F => X"1ac12a031b0129831b4129031b8124031bc120830007851300000793dd8ff0ef",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"1c01011319012d8319412d0319812c8319c12c031a012b831a412b031a812a83",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000008067",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;

--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"0000041300000393000003130000029300000213000001930000011300000093",
        INIT_01 => X"0000081300000793000007130000069300000613000005930000051300000493",
        INIT_02 => X"00000c1300000b9300000b1300000a9300000a13000009930000091300000893",
        INIT_03 => X"0000113700000f9300000f1300000e9300000e1300000d9300000d1300000c93",
        INIT_04 => X"810007b70101041300812623ff0101130000006f001000730080006f6a4000ef",
        INIT_05 => X"000080670101011300c124030000001300e7a02300776713810007b70007a703",
        INIT_06 => X"810007b70007a703810007b7068000ef010104130081242300112623ff010113",
        INIT_07 => X"ff01011300008067010101130081240300c120830000001300e7a02300176713",
        INIT_08 => X"00276713810007b70007a703810007b702c000ef010104130081242300112623",
        INIT_09 => X"00812623ff01011300008067010101130081240300c120830000001300e7a023",
        INIT_0A => X"00c124030000001300e7a023ff877713810007b70007a703810007b701010413",
        INIT_0B => X"00100713000027b7fea426230201041300812e23fe0101130000806701010113",
        INIT_0C => X"0000001300e7a02300700713810007b700e7a02301700713810007b700e7aa23",
        INIT_0D => X"fcb42c23fca42e230301041302812623fd010113000080670201011301c12403",
        INIT_0E => X"00379793fee447830880006ffe0407a31440006ffe040723fcd42823fcc42a23",
        INIT_0F => X"00379793fee4478300e78023fff0071300f707b3fef4478300f70733fdc42703",
        INIT_10 => X"fd44270300379793fee447830007802300f707b3fef4478300f70733fd842703",
        INIT_11 => X"00f70733fd04270300379793fee447830007802300f707b3fef4478300f70733",
        INIT_12 => X"fef44703fef407a300178793fef4478300e78023fff0071300f707b3fef44783",
        INIT_13 => X"fdc4270300379793fee447830880006ffef407a300400793f6e7fae300300793",
        INIT_14 => X"00f70733fd84270300379793fee447830007802300f707b3fef4478300f70733",
        INIT_15 => X"00f70733fd44270300379793fee4478300e78023fff0071300f707b3fef44783",
        INIT_16 => X"fef4478300f70733fd04270300379793fee447830007802300f707b3fef44783",
        INIT_17 => X"00700793fef44703fef407a300178793fef4478300e78023fff0071300f707b3",
        INIT_18 => X"00400793eae7fce300300793fee44703fef4072300178793fee44783f6e7fae3",
        INIT_19 => X"00f70733fdc4270300379793fee447830880006ffe0407a314c0006ffef40723",
        INIT_1A => X"fef4478300f70733fd84270300379793fee447830007802300f707b3fef44783",
        INIT_1B => X"00f707b3fef4478300f70733fd44270300379793fee447830007802300f707b3",
        INIT_1C => X"00f707b3fef4478300f70733fd04270300379793fee4478300e78023fff00713",
        INIT_1D => X"f6e7fae300300793fef44703fef407a300178793fef4478300e78023fff00713",
        INIT_1E => X"fef4478300f70733fdc4270300379793fee447830900006ffef407a300400793",
        INIT_1F => X"fef4478300f70733fd84270300379793fee4478300e7802307f0071300f707b3",
        INIT_20 => X"fef4478300f70733fd44270300379793fee4478300e7802307f0071300f707b3",
        INIT_21 => X"fef4478300f70733fd04270300379793fee4478300e7802307f0071300f707b3",
        INIT_22 => X"00700793fef44703fef407a300178793fef4478300e78023fff0071300f707b3",
        INIT_23 => X"00000013eae7f8e300700793fee44703fef4072300178793fee44783f6e7f6e3",
        INIT_24 => X"fca42e230301041302812623fd010113000080670301011302c1240300000013",
        INIT_25 => X"fdc42783fec4270300078a630017f793fd8427830380006ffe042623fcb42c23",
        INIT_26 => X"fcf42c230017d793fd842783fcf42e2300179793fdc42783fef4262300f707b3",
        INIT_27 => X"fd010113000080670301011302c1240300078513fec42783fc0794e3fd842783",
        INIT_28 => X"fdc42783fef4262300178793fec42783fe042623fca42e230301041302812623",
        INIT_29 => X"0301011302c1240300078513fec42783fe0792e3fdc42783fcf42e234087d793",
        INIT_2A => X"fd442683fcc42a23fcb42e23fca42c230301041302812623fd01011300008067",
        INIT_2B => X"fe068693fec426830980006ffed42623ff868693fe842683fed4242300369693",
        INIT_2C => X"01f0059300169613fdc426830380006f0000079300d65733fdc426030006ca63",
        INIT_2D => X"fec4268300e6e73300c5d733fd842583fec4260300d616b340d586b3fec42683",
        INIT_2E => X"fe442603800006b7fed422230ff6f693fe442683fee4222300d657b3fdc42603",
        INIT_2F => X"00c68823000026b70ff6f613001686930106c683000026b700c680230ff67613",
        INIT_30 => X"02c124030000001300000013f606d4e3fec42683fed42623ff868693fec42683",
        INIT_31 => X"000507930201041300912a2300812c2300112e23fe0101130000806703010113",
        INIT_32 => X"fef4062300070793fef406a300060793fef4072300058793fef407a300068713",
        INIT_33 => X"0007851300500593fee4478300050493e25ff0ef0007851300300593fef44783",
        INIT_34 => X"00050793df9ff0ef0007851300700593fed4478300f484b300050793e11ff0ef",
        INIT_35 => X"03f7f79300f487b300050793de1ff0ef0007851300b00593fec4478300f484b3",
        INIT_36 => X"02812623fd0101130000806702010113014124830181240301c1208300078513",
        INIT_37 => X"00078713fdf44783fcf40f2300070793fcf40fa3000587130005079303010413",
        INIT_38 => X"0301011302c1240300078513fef44783fef407a30ff7f79340f707b3fde44783",
        INIT_39 => X"29512c2329412e232b3120232b2122232a8124232a112623d501011300008067",
        INIT_3A => X"fc0407a32b01041329b1202329a1222329912423298126232971282329612a23",
        INIT_3B => X"e7040693fc042023fcf405a3fff00793fcf40623fff00793fc0406a3fc040723",
        INIT_3C => X"0240006ffa042e23a19ff0ef0007851300070593f3040793ef040713eb040613",
        INIT_3D => X"faf42e2300178793fbc42783da07a023008787b3fd07879300279793fbc42783",
        INIT_3E => X"00e78023000747030007071300002737800007b7fce7dce303f00793fbc42703",
        INIT_3F => X"0007071300002737800007b700e78023001747030007071300002737800007b7",
        INIT_40 => X"000027b700e78023003747030007071300002737800007b700e7802300274703",
        INIT_41 => X"d09ff0efd6c42583d684250300400613d6042623d6f424230047a78300078793",
        INIT_42 => X"d6442583d604250300400613d6042223d6f420230087a78300078793000027b7",
        INIT_43 => X"d584250300100613d4042e23d4f42c2300c7c78300078793000027b7ce5ff0ef",
        INIT_44 => X"0010061300000d9300078d1300d7c78300078793000027b7cc1ff0efd5c42583",
        INIT_45 => X"000027b75d00006ffa040d235f00006ffa040da3c9dff0ef000d8593000d0513",
        INIT_46 => X"fd07879300379793fba44703fbb4478308f71a630040079300c7c70300078793",
        INIT_47 => X"fd07879300379793fba44683fbb4478301879713f607c78300e787b3008787b3",
        INIT_48 => X"00379793fba44683fbb4478300f7673301079793f207c78300d787b3008787b3",
        INIT_49 => X"fba44683fbb4478300f7673300879793ee07c78300d787b3008787b3fd078793",
        INIT_4A => X"06c0006ffcf4222300f767b3ea07c78300d787b3008787b3fd07879300379793",
        INIT_4B => X"01079713f607c78300e787b3008787b3fd07879300379793fba44703fbb44783",
        INIT_4C => X"00879793f207c78300d787b3008787b3fd07879300379793fba44683fbb44783",
        INIT_4D => X"ee07c78300d787b3008787b3fd07879300379793fba44683fbb4478300f76733",
        INIT_4E => X"001787930ff7f793fcb4078300f71e63fc042783fc442703fcf4222300f767b3",
        INIT_4F => X"04f7106303e00793fcb407030007d863fcb4078340c0006ffcf405a30ff7f793",
        INIT_50 => X"ae1ff0ef00078513fa042783faf4222341f7d793faf420230c078793fcb40783",
        INIT_51 => X"fbb44783fcf405a3fff00793b15ff0effa442583fa0425030007861300050793",
        INIT_52 => X"fba44703fbb44783f607c50300e787b3008787b3fd07879300379793fba44703",
        INIT_53 => X"00379793fba44703fbb44783f207c58300e787b3008787b3fd07879300379793",
        INIT_54 => X"fd07879300379793fba44703fbb44783ee07c60300e787b3008787b3fd078793",
        INIT_55 => X"f9f44783f8f40fa300050793b79ff0ef00078693ea07c78300e787b3008787b3",
        INIT_56 => X"0ff7f793f9f4478302f71c63fc442703da07a783008787b3fd07879300279793",
        INIT_57 => X"f70425030007861300050793a0dff0ef00078513f7042783f6042a23f6f42823",
        INIT_58 => X"fc442703008787b3fd07879300279793f9f447832ec0006fa41ff0eff7442583",
        INIT_59 => X"f607c78300e787b3008787b3fd07879300379793fba44703fbb44783dae7a023",
        INIT_5A => X"fba44703fbb44783f8f40f2300050793b8dff0ef0007851300070593fcf44703",
        INIT_5B => X"0007851300070593fce44703f207c78300e787b3008787b3fd07879300379793",
        INIT_5C => X"008787b3fd07879300379793fba44703fbb44783f8f40ea300050793b59ff0ef",
        INIT_5D => X"f8f40e2300050793b25ff0ef0007851300070593fcd44703ee07c78300e787b3",
        INIT_5E => X"ffe00793f9d407030ae7ca6300100793f9e407030cf74063ffe00793f9e40703",
        INIT_5F => X"f9c4070308f74863ffe00793f9c4070308e7ce6300100793f9d407030af74463",
        INIT_60 => X"00e787b3008787b3fd07879300379793fba44703fbb4478308e7c26300100793",
        INIT_61 => X"f9d407830407e7130047979300278793f9e4078306f71063fcc44703ea07c783",
        INIT_62 => X"41f7d793f8f4282300f767b300278793f9c4078300f767330027979300278793",
        INIT_63 => X"f9442583f90425030007861300050793891ff0ef00078513f9042783f8f42a23",
        INIT_64 => X"0ee7c46301f00793f9d407030ef74a63fe000793f9d407031700006f8c5ff0ef",
        INIT_65 => X"40f70733f9d40783f9e407030cf74a63ff80079340f70733f9d40783f9e40703",
        INIT_66 => X"f9c407030af74663ffc0079340f70733f9d40783f9c407030ce7c06300700793",
        INIT_67 => X"fd07879300379793fba44703fbb4478308e7cc630040079340f70733f9d40783",
        INIT_68 => X"0087971302078793f9d4078306f71a63fcc44703ea07c78300e787b3008787b3",
        INIT_69 => X"00f76733004797930087879340f687b3f9d40783f9e4068300f76733000087b7",
        INIT_6A => X"f8f4262341f7d793f8f4242300f767b30087879340f687b3f9d40783f9c40683",
        INIT_6B => X"fc8ff0eff8c42583f88425030007861300050793f94ff0ef00078513f8842783",
        INIT_6C => X"00078913fc44278302f71a630040079300c7c70300078793000027b70740006f",
        INIT_6D => X"f7c42583f784250300500613f7742e23f7642c230ff9eb9300096b1300000993",
        INIT_6E => X"f98420230feaec93000a6c1300000a9300078a13fc4427830300006ff84ff0ef",
        INIT_6F => X"fbb44783fcf42023fc442783f54ff0eff8442583f804250300400613f9942223",
        INIT_70 => X"fbb44783fcf407a3f607c78300e787b3008787b3fd07879300379793fba44703",
        INIT_71 => X"fbb44783fcf40723f207c78300e787b3008787b3fd07879300379793fba44703",
        INIT_72 => X"fbb44783fcf406a3ee07c78300e787b3008787b3fd07879300379793fba44703",
        INIT_73 => X"fba44783fcf40623ea07c78300e787b3008787b3fd07879300379793fba44703",
        INIT_74 => X"faf40da300178793fbb44783a2e7f6e300700793fba44703faf40d2300178793",
        INIT_75 => X"04f7106303e00793fcb407030007d863fcb40783a0e7f6e300700793fbb44703",
        INIT_76 => X"e20ff0ef00078513fb042783faf42a2341f7d793faf428230c078793fcb40783",
        INIT_77 => X"00100713fcf405a3fff00793e54ff0effb442583fb0425030007861300050793",
        INIT_78 => X"00000793e2cff0effac42583fa84250300800613faf42623fae4242300000793",
        INIT_79 => X"29412b0329812a8329c12a032a0129832a4129032a8124032ac1208300078513",
        INIT_7A => X"00000000000080672b01011328012d8328412d0328812c8328c12c0329012b83",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;

--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"0000041300000393000003130000029300000213000001930000011300000093",
        INIT_01 => X"0000081300000793000007130000069300000613000005930000051300000493",
        INIT_02 => X"00000c1300000b9300000b1300000a9300000a13000009930000091300000893",
        INIT_03 => X"0000113700000f9300000f1300000e9300000e1300000d9300000d1300000c93",
        INIT_04 => X"00f720230077e79300072783810007370000006f001000730080006f025000ef",
        INIT_05 => X"00e7a023001767130007a70300e7a023ff8777130007a703810007b700008067",
        INIT_06 => X"00e7a023002767130007a70300e7a023ff8777130007a703810007b700008067",
        INIT_07 => X"00100713000027b70000806700f72023ff87f793000727838100073700008067",
        INIT_08 => X"007587930000806700e7a0230070071300e7a02301700713810007b700e7a823",
        INIT_09 => X"0018381340d7073300f8381300f33313007507930076071340c7883340d78333",
        INIT_0A => X"0067773300f8b89340c78833001737130103733300f737130013331340b788b3",
        INIT_0B => X"01177733ff0101130018371300f7b79300e8f8b340d787b300f838130018b893",
        INIT_0C => X"00f5e7b300d667b32007806300e7f7b30121222300912423008126230017b793",
        INIT_0D => X"00f5a2230005a0230005222300f52023fff007931e0796630037f79300f567b3",
        INIT_0E => X"00f5a6230005a4230005262300f5242300f6a22300f6a0230006222300062023",
        INIT_0F => X"00f5aa230005a82300052a2300f5282300f6a62300f6a4230006262300062423",
        INIT_10 => X"00f5ae230005ac2300052e2300f52c2300f6aa2300f6a82300062a2300062823",
        INIT_11 => X"0285889302068e1302060e930205831300f6ae2300f6ac2300062e2300062c23",
        INIT_12 => X"0285071302050f13011e343301f333b3011eb933010337b302868f9302860813",
        INIT_13 => X"0127e7b30083e3b30013b393001939130017b79301feb4b3010e32b300143413",
        INIT_14 => X"0018b89300eeb3b30092e2b30077f7b3011f38b30014b4930012b29300e33433",
        INIT_15 => X"01ff3fb300ee37330013b293001838130088e8b30057f7b3010f383300143413",
        INIT_16 => X"2c07806300e7f7b301f767330107f7b3001fbf9300173713005868330117f7b3",
        INIT_17 => X"02052023f7f787937f7f87b72a0f1663003f7f13006f6f3301c3633301de6e33",
        INIT_18 => X"02e6a22302e6a02302f6222302e62023fff0071302f5a2230205a02302f52223",
        INIT_19 => X"02e6a62302e6a42302f6262302e6242302f5a6230205a42302f5262302052423",
        INIT_1A => X"02e6aa2302e6a82302f62a2302e6282302f5aa230205a82302f52a2302052823",
        INIT_1B => X"02e6ae2302e6ac2302f62e2302e62c2302f5ae230205ac2302f52e2302052c23",
        INIT_1C => X"0005802300f50023fff007930000806701010113004129030081248300c12403",
        INIT_1D => X"0005812300f5012300f680a3000600a3000580a300f500a300f6802300060023",
        INIT_1E => X"00f582230005022300f681a3000601a3000581a300f501a300f6812300060123",
        INIT_1F => X"00f583230005032300f682a3000602a300f582a3000502a300f6822300060223",
        INIT_20 => X"0005842300f5042300f683a3000603a300f583a3000503a300f6832300060323",
        INIT_21 => X"0005852300f5052300f684a3000604a3000584a300f504a300f6842300060423",
        INIT_22 => X"00f586230005062300f685a3000605a3000585a300f505a300f6852300060523",
        INIT_23 => X"00f587230005072300f686a3000606a300f586a3000506a300f6862300060623",
        INIT_24 => X"0005882300f5082300f687a3000607a300f587a3000507a300f6872300060723",
        INIT_25 => X"0005892300f5092300f688a3000608a3000588a300f508a300f6882300060823",
        INIT_26 => X"00f58a2300050a2300f689a3000609a3000589a300f509a300f6892300060923",
        INIT_27 => X"00f58b2300050b2300f68aa300060aa300f58aa300050aa300f68a2300060a23",
        INIT_28 => X"00058c2300f50c2300f68ba300060ba300f58ba300050ba300f68b2300060b23",
        INIT_29 => X"00058d2300f50d2300f68ca300060ca300058ca300f50ca300f68c2300060c23",
        INIT_2A => X"00f58e2300050e2300f68da300060da300058da300f50da300f68d2300060d23",
        INIT_2B => X"00f58f2300050f2300f68ea300060ea300f58ea300050ea300f68e2300060e23",
        INIT_2C => X"02050023c99ff06f00f68fa300060fa300f58fa300050fa300f68f2300060f23",
        INIT_2D => X"02f680a302f600a3020580a3020500a302f6802302f6002302058023fff00793",
        INIT_2E => X"07f0071302f601a3020581a3020501a302f6812302f601230205812302050123",
        INIT_2F => X"02e602a302e582a302e502a302f6822302e6022302e5822302e5022302f681a3",
        INIT_30 => X"02e603a302e583a302e503a302f6832302e6032302e5832302e5032302f682a3",
        INIT_31 => X"02f604a3020584a3020504a302f6842302f60423020584230205042302f683a3",
        INIT_32 => X"02f605a3020585a3020505a302f6852302f60523020585230205052302f684a3",
        INIT_33 => X"02e606a302e586a302e506a302f6862302e6062302e5862302e5062302f685a3",
        INIT_34 => X"02e607a302e587a302e507a302f6872302e6072302e5872302e5072302f686a3",
        INIT_35 => X"02f608a3020588a3020508a302f6882302f60823020588230205082302f687a3",
        INIT_36 => X"02f609a3020589a3020509a302f6892302f60923020589230205092302f688a3",
        INIT_37 => X"02e60aa302e58aa302e50aa302f68a2302e60a2302e58a2302e50a2302f689a3",
        INIT_38 => X"02e60ba302e58ba302e50ba302f68b2302e60b2302e58b2302e50b2302f68aa3",
        INIT_39 => X"02f60ca302058ca302050ca302f68c2302f60c2302058c2302050c2302f68ba3",
        INIT_3A => X"02f60da302058da302050da302f68d2302f60d2302058d2302050d2302f68ca3",
        INIT_3B => X"02e60ea302e58ea302e50ea302f68e2302e60e2302e58e2302e50e2302f68da3",
        INIT_3C => X"00c1240302e58fa302e50fa302f68f2302e60f2302e58f2302e50f2302f68ea3",
        INIT_3D => X"00000513000507930000806701010113004129030081248302f68fa302e60fa3",
        INIT_3E => X"00008067fe0596e30017979300f50533000704630015d5930015f71302058063",
        INIT_3F => X"0036161300008067fe079ce3001505134087d793000005130005079300008067",
        INIT_40 => X"00c5573340c307b3800008b701f0031300159e130000283704064663ff860613",
        INIT_41 => X"0148478300e880230ff7771300d5d7330006c46300e7e733fe06069300fe17b3",
        INIT_42 => X"00d787b300c787b30016979300008067fc0656e300f80a2300178793ff860613",
        INIT_43 => X"0025959300d787b30036969300c787b30026161300e787b300b787b300161713",
        INIT_44 => X"0ff5751340b505330000806703f5751300e7853300a7073300b787b300151713",
        INIT_45 => X"24812423241126230101051305010593090106130d010693db01011300008067",
        INIT_46 => X"23812423237126232361282323512a2323412c2323312e232521202324912223",
        INIT_47 => X"004787930007a0232101071311010793831ff0ef21b12e2323a1202323912223",
        INIT_48 => X"00e78023002a4603001a4583800007b7000a4703000a0a1300002a37fef71ce3",
        INIT_49 => X"000025b700d780230187569300d7802300c7802300b78023003a4683004a2703",
        INIT_4A => X"008756930145c60300d7802300c58a23001606130ff6f693010756930145c603",
        INIT_4B => X"00160613008a27030ff776930145c60300d7802300c58a23001606130ff6f693",
        INIT_4C => X"00a7802300d58a230016869301075613018755130145c68300d7802300c58a23",
        INIT_4D => X"0ff6f6930145c60300c7802300a58a2300150513008756930ff676130145c503",
        INIT_4E => X"0016869305010413090109130145c68300d7802300c58a23001606130ff77713",
        INIT_4F => X"00c7802300e58a230017071300da468300ca46030145c70300e7802300d58a23",
        INIT_50 => X"000007930145c70300d7802300e58a23001707130d010b9301810b130145c703",
        INIT_51 => X"0000069300000313000409130ff00c930009071300e58a2300170713fff00393",
        INIT_52 => X"00ca4783000786130007041301f00d9380000eb700300d1300400a9300000813",
        INIT_53 => X"000fc883000e440301712623012122230081242300090f93ff8b0e1300040293",
        INIT_54 => X"00e7e7b3008897130104179317578e630080099303f00c13000b8f130002c503",
        INIT_55 => X"002514930126063300a4063300289713000f49033203de6318c7846300a7e7b3",
        INIT_56 => X"03f77713009707330177073300c484b30016149300391b930097073301170733",
        INIT_57 => X"4104083320f48e630ff77713f006248300960633200606130101049300271613",
        INIT_58 => X"0ff6f7130ff375130ff7761301881813f0f620234065033340d886b300280713",
        INIT_59 => X"32c6c463ffe0061320cd6063418353134186d693418858130186969301831313",
        INIT_5A => X"ff80069340e8083300d66e6303f006130ff6f6930207069342d8de6300100893",
        INIT_5B => X"00ee80230187d7131557006300ca47031ed55c63ffc0069340e3053300d84863",
        INIT_5C => X"0087d7130145c68300ee802300d58a23001686930ff777130107d7130145c683",
        INIT_5D => X"00d58a23001686930ff7f7130145c68300ee802300d58a23001686930ff77713",
        INIT_5E => X"001e0e1300e58a23001707130002c303000fc683000e48030145c70300ee8023",
        INIT_5F => X"000e440300ca47830007861307cb0663001f0f1300128293001f8f93000f4c83",
        INIT_60 => X"00e7e7b30097e7b30108949301841793000f4703e95796e30002c503000fc883",
        INIT_61 => X"4183d393000f4c83001e0e130183939300138393e8c790e300e7e7b300851713",
        INIT_62 => X"00412903f9cb1ee3001f0f1300128293001f8f93000408130008869300050313",
        INIT_63 => X"dd271ee3008b8b9300840413008b0b13090107130089091300c12b8300812403",
        INIT_64 => X"00179513fd87069341f3d79300371713001707134083d7130c0383932203cc63",
        INIT_65 => X"0145c60300ee8023fff007131d80006f1e06d86300d7d7b300800613ff870713",
        INIT_66 => X"0087d7130ff6f6930145c60300ee802300c58a23001606130107d6930187d713",
        INIT_67 => X"00c58a23001606130ff7f6930ff777130145c60300de802300c58a2300160613",
        INIT_68 => X"000e48030145c70300ee80230006871300e58a23001707130145c70300ee8023",
        INIT_69 => X"e2ec6ae30ff7771302070713eadff06f00e58a230002c30300170713000fc683",
        INIT_6A => X"ffc0069340e30533e106cee300700693e2d842e3ff80069340d8083300068713",
        INIT_6B => X"00d7673300871713004816930207071300880813e19914e3e0aac6e3e0d548e3",
        INIT_6C => X"0080006f008008130080069341f7589300d7673300a76733000086b700850513",
        INIT_6D => X"0ff6761300c566330065153300d756330018951340d3033301f0031300000693",
        INIT_6E => X"0002c303000fc683000e4803fd0688e300c58a23001606130145c60300ce8023",
        INIT_6F => X"00171513fd86089341f3d71300361613001606134083d6130c038393dfdff06f",
        INIT_70 => X"00e58a23001707130145c70300ee80230ff777130208c06301175733ff860613",
        INIT_71 => X"00ee80230ff7771300e8e73300c3d733011518b340cd88b30000061303361863",
        INIT_72 => X"fff00393000fc8830002c503000e4403fd360ce300e58a23001707130145c703",
        INIT_73 => X"cf06cae30070069340d8083300068713d0ec62e30ff7771302070713c4dff06f",
        INIT_74 => X"0ff7f79300f6e7b300e3d7b300d516b340e686b301f0069300000713ed9ff06f",
        INIT_75 => X"00078023800007b7fcc708e300f58a23001787930145c78300f68023800006b7",
        INIT_76 => X"00e58a23001707130145c7030007802300e58a2300170713000005130145c703",
        INIT_77 => X"00e58a23001707130145c7030007802300e58a23001707130145c70300078023",
        INIT_78 => X"00e58a23001707130145c7030007802300e58a23001707130145c70300078023",
        INIT_79 => X"248124030145c78300e780230010071300e58a23001707130145c70300078023",
        INIT_7A => X"23012b0323412a8323812a0323c1298324012903244124830017879324c12083",
        INIT_7B => X"000080672501011321c12d8322012d0322412c8322812c0322c12b8300f58a23",
        INIT_7C => X"00068713dd1ff06fbcaacee340d808330006871340d505330268da6300c34e63",
        INIT_7D => X"00280713bb991ce3db9ff06fbd9910e3bcd542e340e80833ffc0069340d30533",
        INIT_7E => X"0ff7771304076713006767330023031300d76733004717130026969300268693",
        INIT_7F => X"0000000000000000000000000000000000000000d31ff06f00e68023800006b7",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;

--------------------------------------------------------------------------------
-- KU Leuven - ESAT/COSIC - Emerging technologies, Systems & Security
--------------------------------------------------------------------------------
-- Module Name:     two_k_bram_imem - Behavioural
-- Project Name:    two_k_bram_imem
-- Description:     
--
-- Revision     Date       Author     Comments
-- v0.1         20250204   VlJo       Initial version
--
--------------------------------------------------------------------------------
library IEEE;
    use IEEE.STD_LOGIC_1164.ALL;
    -- use IEEE.NUMERIC_STD.ALL;

Library UNISIM;
    use UNISIM.vcomponents.all;

entity two_k_bram_imem is
    port(
        clock : in STD_LOGIC;

        init_data_in : in STD_LOGIC_VECTOR(31 downto 0);
        init_write_enable : in STD_LOGIC;
        init_address : in STD_LOGIC_VECTOR(10 downto 0);

        data_in : in STD_LOGIC_VECTOR(31 downto 0);
        write_enable : in STD_LOGIC;
        address : in STD_LOGIC_VECTOR(10 downto 0);
        data_out : out STD_LOGIC_VECTOR(31 downto 0)
    );
end entity two_k_bram_imem;

architecture Behavioural of two_k_bram_imem is

    -- (DE-)LOCALISING IN/OUTPUTS
    signal clock_i : STD_LOGIC;
    signal init_data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal init_write_enable_i : STD_LOGIC;
    signal init_address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_in_i : STD_LOGIC_VECTOR(31 downto 0);
    signal write_enable_i : STD_LOGIC;
    signal address_i : STD_LOGIC_VECTOR(10 downto 0);
    signal data_out_o : STD_LOGIC_VECTOR(31 downto 0);

    constant C_NULL : STD_LOGIC_VECTOR(31 downto 0) := x"00000000";
    constant C_ONES : STD_LOGIC_VECTOR(31 downto 0) := x"FFFFFFFF";

    signal init_address_00, init_address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal init_write_enable_00, init_write_enable_01 : STD_LOGIC;
    signal init_write_enable_00_vec, init_write_enable_01_vec : STD_LOGIC_VECTOR(3 downto 0);

    signal address_00, address_01 : STD_LOGIC_VECTOR(15 downto 0);
    signal write_enable_00, write_enable_01 : STD_LOGIC;
    signal write_enable_00_vec, write_enable_01_vec : STD_LOGIC_VECTOR(7 downto 0);
    signal data_out_00, data_out_01 : STD_LOGIC_VECTOR(31 downto 0);


begin

    -------------------------------------------------------------------------------
    -- (DE-)LOCALISING IN/OUTPUTS
    -------------------------------------------------------------------------------
    clock_i <= clock;
    init_data_in_i <= init_data_in;
    init_write_enable_i <= init_write_enable;
    init_address_i <= init_address;

    data_in_i <= data_in;
    write_enable_i <= write_enable;
    address_i <= address;
    data_out <= data_out_o;


    init_address_00 <= "0" & init_address_i(9 downto 0) & "00000";
    init_address_01 <= "0" & init_address_i(9 downto 0) & "00000";
    init_write_enable_00 <= init_write_enable_i and not(init_address(10));
    init_write_enable_01 <= init_write_enable_i and init_address(10);    
    init_write_enable_00_vec <= (others => init_write_enable_00);
    init_write_enable_01_vec <= (others => init_write_enable_01);
    
    address_00 <= "0" & address_i(9 downto 0) & "00000";
    address_01 <= "0" & address_i(9 downto 0) & "00000";
    write_enable_00 <= write_enable_i and not(address_i(10));
    write_enable_01 <= write_enable_i and address_i(10);
    write_enable_00_vec <= (others => write_enable_00);
    write_enable_01_vec <= (others => write_enable_01);
    data_out_o <= data_out_00 when address_i(10) = '0' else data_out_01;
    

    -------------------------------------------------------------------------------
    -- BRAM PRIMITIVES
    -------------------------------------------------------------------------------
    RAMB36E1_inst00 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"004124230031222300112023340111730000001300000013000000131140006f",
        INIT_01 => X"02c1242302b1222302a1202300912e2300812c2300712a230061282300512623",
        INIT_02 => X"05412423053122230521202303112e2303012c2302f12a2302e1282302d12623",
        INIT_03 => X"07c1242307b1222307a1202305912e2305812c2305712a230561282305512623",
        INIT_04 => X"008122030041218300012083278000ef3420357307f12a2307e1282307d12623",
        INIT_05 => X"02812603024125830201250301c1248301812403014123830101230300c12283",
        INIT_06 => X"04812a03044129830401290303c1288303812803034127830301270302c12683",
        INIT_07 => X"06812e0306412d8306012d0305c12c8305812c0305412b8305012b0304c12a83",
        INIT_08 => X"000001930000011300000093302000733401117307412f8307012f0306c12e83",
        INIT_09 => X"0000059300000513000004930000041300000393000003130000029300000213",
        INIT_0A => X"0000099300000913000008930000081300000793000007130000069300000613",
        INIT_0B => X"00000d9300000d1300000c9300000c1300000b9300000b1300000a9300000a13",
        INIT_0C => X"eef18193deadc1b7fe0101130000113700000f9300000f1300000e9300000e13",
        INIT_0D => X"3004507330511073e60101130000011734011073000101130000113700018213",
        INIT_0E => X"00112023ff4101130540006f708000ef00100073710000ef30411073fff00113",
        INIT_0F => X"0005853300029663fff50293000583330280006f000514630061242300512223",
        INIT_10 => X"00812303004122830001208300030533fe029ce3fff2829300b303330140006f",
        INIT_11 => X"810007b70101041300812623ff0101130000006f0000006f0000806700c10113",
        INIT_12 => X"000080670101011300c124030000001300e7a02300776713810007b70007a703",
        INIT_13 => X"810007b70007a703810007b7068000ef010104130081242300112623ff010113",
        INIT_14 => X"ff01011300008067010101130081240300c120830000001300e7a02300176713",
        INIT_15 => X"00276713810007b70007a703810007b702c000ef010104130081242300112623",
        INIT_16 => X"00812623ff01011300008067010101130081240300c120830000001300e7a023",
        INIT_17 => X"00c124030000001300e7a023ff877713810007b70007a703810007b701010413",
        INIT_18 => X"00100713000027b7fea426230201041300812e23fe0101130000806701010113",
        INIT_19 => X"0000001300e7a02300700713810007b700e7a02301700713810007b700e7aa23",
        INIT_1A => X"fcb42c23fca42e230301041302812623fd010113000080670201011301c12403",
        INIT_1B => X"00379793fee447830880006ffe0407a31440006ffe040723fcd42823fcc42a23",
        INIT_1C => X"00379793fee4478300e78023fff0071300f707b3fef4478300f70733fdc42703",
        INIT_1D => X"fd44270300379793fee447830007802300f707b3fef4478300f70733fd842703",
        INIT_1E => X"00f70733fd04270300379793fee447830007802300f707b3fef4478300f70733",
        INIT_1F => X"fef44703fef407a300178793fef4478300e78023fff0071300f707b3fef44783",
        INIT_20 => X"fdc4270300379793fee447830880006ffef407a300400793f6e7fae300300793",
        INIT_21 => X"00f70733fd84270300379793fee447830007802300f707b3fef4478300f70733",
        INIT_22 => X"00f70733fd44270300379793fee4478300e78023fff0071300f707b3fef44783",
        INIT_23 => X"fef4478300f70733fd04270300379793fee447830007802300f707b3fef44783",
        INIT_24 => X"00700793fef44703fef407a300178793fef4478300e78023fff0071300f707b3",
        INIT_25 => X"00400793eae7fce300300793fee44703fef4072300178793fee44783f6e7fae3",
        INIT_26 => X"00f70733fdc4270300379793fee447830880006ffe0407a314c0006ffef40723",
        INIT_27 => X"fef4478300f70733fd84270300379793fee447830007802300f707b3fef44783",
        INIT_28 => X"00f707b3fef4478300f70733fd44270300379793fee447830007802300f707b3",
        INIT_29 => X"00f707b3fef4478300f70733fd04270300379793fee4478300e78023fff00713",
        INIT_2A => X"f6e7fae300300793fef44703fef407a300178793fef4478300e78023fff00713",
        INIT_2B => X"fef4478300f70733fdc4270300379793fee447830900006ffef407a300400793",
        INIT_2C => X"fef4478300f70733fd84270300379793fee4478300e7802307f0071300f707b3",
        INIT_2D => X"fef4478300f70733fd44270300379793fee4478300e7802307f0071300f707b3",
        INIT_2E => X"fef4478300f70733fd04270300379793fee4478300e7802307f0071300f707b3",
        INIT_2F => X"00700793fef44703fef407a300178793fef4478300e78023fff0071300f707b3",
        INIT_30 => X"00000013eae7f8e300700793fee44703fef4072300178793fee44783f6e7f6e3",
        INIT_31 => X"fca42e230301041302812623fd010113000080670301011302c1240300000013",
        INIT_32 => X"fdc42783fec4270300078a630017f793fd8427830380006ffe042623fcb42c23",
        INIT_33 => X"fcf42c230017d793fd842783fcf42e2300179793fdc42783fef4262300f707b3",
        INIT_34 => X"fd010113000080670301011302c1240300078513fec42783fc0794e3fd842783",
        INIT_35 => X"fdc42783fef4262300178793fec42783fe042623fca42e230301041302812623",
        INIT_36 => X"0301011302c1240300078513fec42783fe0792e3fdc42783fcf42e234087d793",
        INIT_37 => X"fd442683fcc42a23fcb42e23fca42c230301041302812623fd01011300008067",
        INIT_38 => X"fe068693fec426830ac0006ffed42623ff868693fe842683fed4242300369693",
        INIT_39 => X"01f0059300169613fdc426830380006f0000079300d65733fdc426030006ca63",
        INIT_3A => X"fec4268300e6e73300c5d733fd842583fec4260300d616b340d586b3fec42683",
        INIT_3B => X"0106c683000026b7fed422230ff6f693fe442683fee4222300d657b3fdc42603",
        INIT_3C => X"000026b700d600230ff6f693fe4426830006861300d606b3800006b700068613",
        INIT_3D => X"fed42623ff868693fec4268300c68823000026b70ff6f613001686930106c683",
        INIT_3E => X"fe010113000080670301011302c124030000001300000013f406dae3fec42683",
        INIT_3F => X"00058793fef407a300068713000507930201041300912a2300812c2300112e23",
        INIT_40 => X"0007851300300593fef44783fef4062300070793fef406a300060793fef40723",
        INIT_41 => X"00f484b300050793dfdff0ef0007851300500593fee4478300050493e11ff0ef",
        INIT_42 => X"00b00593fec4478300f484b300050793de5ff0ef0007851300700593fed44783",
        INIT_43 => X"0181240301c120830007851303f7f79300f487b300050793dcdff0ef00078513",
        INIT_44 => X"00058713000507930301041302812623fd010113000080670201011301412483",
        INIT_45 => X"0ff7f79340f707b3fde4478300078713fdf44783fcf40f2300070793fcf40fa3",
        INIT_46 => X"2a112623d5010113000080670301011302c1240300078513fef44783fef407a3",
        INIT_47 => X"298126232971282329612a2329512c2329412e232b3120232b2122232a812423",
        INIT_48 => X"fff00793fc0406a3fc040723fc0407a32b01041329b1202329a1222329912423",
        INIT_49 => X"f3040793ef040713eb040613e7040693fc042023fcf405a3fff00793fcf40623",
        INIT_4A => X"fd07879300279793fbf447830240006ffa040fa3a05ff0ef0007851300070593",
        INIT_4B => X"fce7fce303f00793fbf44703faf40fa300178793fbf44783da07a023008787b3",
        INIT_4C => X"00e6873380000737000706930107470300002737fbe447830580006ffa040f23",
        INIT_4D => X"0107c783000027b700f680230007c78300f707b3000707130000273700070693",
        INIT_4E => X"fbe44703faf40f2300178793fbe4478300e78823000027b70ff7f71300178793",
        INIT_4F => X"00400613d6042623d6f424230047a78300078793000027b7fae7f2e300300793",
        INIT_50 => X"d6042223d6f420230087a78300078793000027b7cddff0efd6c42583d6842503",
        INIT_51 => X"d4f42c2300c7c78300078793000027b7cb9ff0efd6442583d604250300400613",
        INIT_52 => X"00d7c78300078793000027b7c95ff0efd5c42583d584250300100613d4042e23",
        INIT_53 => X"5f00006ffa040ea3c71ff0ef000d8593000d05130010061300000d9300078d13",
        INIT_54 => X"fbd4478308f71a630040079300c7c70300078793000027b75d00006ffa040e23",
        INIT_55 => X"fbd4478301879713f607c78300e787b3008787b3fd07879300379793fbc44703",
        INIT_56 => X"00f7673301079793f207c78300d787b3008787b3fd07879300379793fbc44683",
        INIT_57 => X"00879793ee07c78300d787b3008787b3fd07879300379793fbc44683fbd44783",
        INIT_58 => X"ea07c78300d787b3008787b3fd07879300379793fbc44683fbd4478300f76733",
        INIT_59 => X"008787b3fd07879300379793fbc44703fbd4478306c0006ffcf4222300f767b3",
        INIT_5A => X"008787b3fd07879300379793fbc44683fbd4478301079713f607c78300e787b3",
        INIT_5B => X"fd07879300379793fbc44683fbd4478300f7673300879793f207c78300d787b3",
        INIT_5C => X"00f71e63fc042783fc442703fcf4222300f767b3ee07c78300d787b3008787b3",
        INIT_5D => X"0007d863fcb4078340c0006ffcf405a30ff7f793001787930ff7f793fcb40783",
        INIT_5E => X"faf4222341f7d793faf420230c078793fcb4078304f7106303e00793fcb40703",
        INIT_5F => X"ae9ff0effa442583fa0425030007861300050793ab5ff0ef00078513fa042783",
        INIT_60 => X"00e787b3008787b3fd07879300379793fbc44703fbd44783fcf405a3fff00793",
        INIT_61 => X"f207c58300e787b3008787b3fd07879300379793fbc44703fbd44783f607c503",
        INIT_62 => X"fbd44783ee07c60300e787b3008787b3fd07879300379793fbc44703fbd44783",
        INIT_63 => X"b61ff0ef00078693ea07c78300e787b3008787b3fd07879300379793fbc44703",
        INIT_64 => X"fc442703da07a783008787b3fd07879300279793f9f44783f8f40fa300050793",
        INIT_65 => X"9e1ff0ef00078513f7042783f6042a23f6f428230ff7f793f9f4478302f71c63",
        INIT_66 => X"00279793f9f447832ec0006fa15ff0eff7442583f70425030007861300050793",
        INIT_67 => X"fd07879300379793fbc44703fbd44783dae7a023fc442703008787b3fd078793",
        INIT_68 => X"00050793b75ff0ef0007851300070593fcf44703f607c78300e787b3008787b3",
        INIT_69 => X"f207c78300e787b3008787b3fd07879300379793fbc44703fbd44783f8f40f23",
        INIT_6A => X"fbc44703fbd44783f8f40ea300050793b41ff0ef0007851300070593fce44703",
        INIT_6B => X"0007851300070593fcd44703ee07c78300e787b3008787b3fd07879300379793",
        INIT_6C => X"00100793f9e407030cf74063ffe00793f9e40703f8f40e2300050793b0dff0ef",
        INIT_6D => X"f9c4070308e7ce6300100793f9d407030af74463ffe00793f9d407030ae7ca63",
        INIT_6E => X"00379793fbc44703fbd4478308e7c26300100793f9c4070308f74863ffe00793",
        INIT_6F => X"00278793f9e4078306f71063fcc44703ea07c78300e787b3008787b3fd078793",
        INIT_70 => X"00278793f9c4078300f767330027979300278793f9d407830407e71300479793",
        INIT_71 => X"00050793865ff0ef00078513f9042783f8f42a2341f7d793f8f4282300f767b3",
        INIT_72 => X"0ef74a63fe000793f9d407031700006f899ff0eff9442583f904250300078613",
        INIT_73 => X"0cf74a63ff80079340f70733f9d40783f9e407030ee7c46301f00793f9d40703",
        INIT_74 => X"40f70733f9d40783f9c407030ce7c0630070079340f70733f9d40783f9e40703",
        INIT_75 => X"fbd4478308e7cc630040079340f70733f9d40783f9c407030af74663ffc00793",
        INIT_76 => X"06f71a63fcc44703ea07c78300e787b3008787b3fd07879300379793fbc44703",
        INIT_77 => X"40f687b3f9d40783f9e4068300f76733000087b70087971302078793f9d40783",
        INIT_78 => X"00f767b30087879340f687b3f9d40783f9c4068300f767330047979300878793",
        INIT_79 => X"0007861300050793f68ff0ef00078513f8842783f8f4262341f7d793f8f42423",
        INIT_7A => X"0040079300c7c70300078793000027b70740006ff9cff0eff8c42583f8842503",
        INIT_7B => X"f7742e23f7642c230ff9eb9300096b130000099300078913fc44278302f71a63",
        INIT_7C => X"00000a9300078a13fc4427830300006ff58ff0eff7c42583f784250300500613",
        INIT_7D => X"f28ff0eff8442583f804250300400613f9942223f98420230feaec93000a6c13",
        INIT_7E => X"00e787b3008787b3fd07879300379793fbc44703fbd44783fcf42023fc442783",
        INIT_7F => X"00e787b3008787b3fd07879300379793fbc44703fbd44783fcf407a3f607c783",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_00,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_00,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_00_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_00,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_00_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

    RAMB36E1_inst01 : RAMB36E1
    generic map (
        RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
        SIM_COLLISION_CHECK => "ALL",
        DOA_REG => 0,
        DOB_REG => 0,
        EN_ECC_READ => FALSE,
        EN_ECC_WRITE => FALSE,
        -- INIT_00 to INIT_7F: Initial contents of the data memory array
        INIT_00 => X"00e787b3008787b3fd07879300379793fbc44703fbd44783fcf40723f207c783",
        INIT_01 => X"00e787b3008787b3fd07879300379793fbc44703fbd44783fcf406a3ee07c783",
        INIT_02 => X"a2e7f6e300700793fbc44703faf40e2300178793fbc44783fcf40623ea07c783",
        INIT_03 => X"0007d863fcb40783a0e7f6e300700793fbd44703faf40ea300178793fbd44783",
        INIT_04 => X"faf42a2341f7d793faf428230c078793fcb4078304f7106303e00793fcb40703",
        INIT_05 => X"e28ff0effb442583fb0425030007861300050793df4ff0ef00078513fb042783",
        INIT_06 => X"fa84250300800613faf42623fae424230000079300100713fcf405a3fff00793",
        INIT_07 => X"2a0129832a4129032a8124032ac120830007851300000793e00ff0effac42583",
        INIT_08 => X"28012d8328412d0328812c8328c12c0329012b8329412b0329812a8329c12a03",
        INIT_09 => X"000000000000000000000000000000000000000000000000000080672b010113",
        INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",
        INIT_A => X"000000000",
        INIT_B => X"000000000",
        INIT_FILE => "NONE",
        RAM_MODE => "TDP", -- RAM Mode: "SDP" or "TDP" 
        RAM_EXTENSION_A => "NONE", -- RAM_EXTENSION_A, RAM_EXTENSION_B: Selects cascade mode ("UPPER", "LOWER", or "NONE")
        RAM_EXTENSION_B => "NONE",
        READ_WIDTH_A => 36, -- 0-72
        READ_WIDTH_B => 36, -- 0-36
        WRITE_WIDTH_A => 36, -- 0-36
        WRITE_WIDTH_B => 36, -- 0-72
        RSTREG_PRIORITY_A => "RSTREG", ---- RSTREG_PRIORITY_A, RSTREG_PRIORITY_B: Reset or enable priority ("RSTREG" or "REGCE")
        RSTREG_PRIORITY_B => "RSTREG",
        SRVAL_A => X"000000000", -- SRVAL_A, SRVAL_B: Set/reset value for output
        SRVAL_B => X"000000000",
        SIM_DEVICE => "7SERIES",
        WRITE_MODE_A => "WRITE_FIRST",  -- WriteMode: Value on output upon a write ("WRITE_FIRST", "READ_FIRST", or "NO_CHANGE")
        WRITE_MODE_B => "WRITE_FIRST" 
    )
   port map (
        CASCADEOUTA => open,
        CASCADEOUTB => open,
        DBITERR => open,
        ECCPARITY => open,
        RDADDRECC => open,
        SBITERR => open,
        DOADO => open,
        DOPADOP => open,
        DOBDO => data_out_01,
        DOPBDOP => open,
        CASCADEINA => C_NULL(0),
        CASCADEINB => C_NULL(0),
        INJECTDBITERR => C_NULL(0),
        INJECTSBITERR => C_NULL(0),
        ADDRARDADDR => init_address_01,
        CLKARDCLK => clock_i,
        ENARDEN => C_NULL(0),
        REGCEAREGCE => C_NULL(0),
        RSTRAMARSTRAM => C_NULL(0),
        RSTREGARSTREG => C_NULL(0),
        WEA => init_write_enable_01_vec,
        DIADI => init_data_in_i,
        DIPADIP => C_NULL(3 downto 0),
        ADDRBWRADDR => address_01,
        CLKBWRCLK => clock_i,
        ENBWREN => C_ONES(0),
        REGCEB => C_NULL(0),
        RSTRAMB => C_NULL(0),
        RSTREGB => C_NULL(0),
        WEBWE => write_enable_01_vec,
        DIBDI => data_in_i,
        DIPBDIP => C_NULL(3 downto 0)
    );

end Behavioural;
